magic
tech sky130A
magscale 1 2
timestamp 1715771064
<< metal1 >>
rect 18750 16650 19050 16656
rect 19050 16350 19942 16650
rect 18750 16344 19050 16350
rect 30532 8340 31140 8500
rect 30532 8160 31462 8340
rect 30532 8040 31140 8160
rect 31282 8120 31462 8160
rect 31276 7940 31282 8120
rect 31462 7940 31468 8120
<< via1 >>
rect 18750 16350 19050 16650
rect 31282 7940 31462 8120
<< metal2 >>
rect 18055 16650 18345 16654
rect 18050 16645 18750 16650
rect 18050 16355 18055 16645
rect 18345 16355 18750 16645
rect 18050 16350 18750 16355
rect 19050 16350 19056 16650
rect 18055 16346 18345 16350
rect 13355 9050 13645 9054
rect 13350 9045 19942 9050
rect 13350 8755 13355 9045
rect 13645 8755 19942 9045
rect 13350 8750 19942 8755
rect 13355 8746 13645 8750
rect 31282 8120 31462 8126
rect 31282 6985 31462 7940
rect 31278 6815 31287 6985
rect 31457 6815 31466 6985
rect 31282 6810 31462 6815
<< via2 >>
rect 18055 16355 18345 16645
rect 13355 8755 13645 9045
rect 31287 6815 31457 6985
<< metal3 >>
rect 17451 16650 17749 16655
rect 17450 16649 18350 16650
rect 17450 16351 17451 16649
rect 17749 16645 18350 16649
rect 17749 16355 18055 16645
rect 18345 16355 18350 16645
rect 17749 16351 18350 16355
rect 17450 16350 18350 16351
rect 17451 16345 17749 16350
rect 5651 9050 5949 9055
rect 5650 9049 13650 9050
rect 5650 8751 5651 9049
rect 5949 9045 13650 9049
rect 5949 8755 13355 9045
rect 13645 8755 13650 9045
rect 5949 8751 13650 8755
rect 5650 8750 13650 8751
rect 5651 8745 5949 8750
rect 31282 6985 31462 6990
rect 31282 6815 31287 6985
rect 31457 6815 31462 6985
rect 31282 1729 31462 6815
rect 31277 1551 31283 1729
rect 31461 1551 31467 1729
rect 31282 1550 31462 1551
<< via3 >>
rect 17451 16351 17749 16649
rect 5651 8751 5949 9049
rect 31283 1551 31461 1729
<< metal4 >>
rect 798 44760 858 45152
rect 1534 44760 1594 45152
rect 2270 44760 2330 45152
rect 3006 44760 3066 45152
rect 3742 44760 3802 45152
rect 4478 44760 4538 45152
rect 5214 44760 5274 45152
rect 5950 44760 6010 45152
rect 6686 44760 6746 45152
rect 7422 44760 7482 45152
rect 8158 44760 8218 45152
rect 8894 44760 8954 45152
rect 9630 44760 9690 45152
rect 10366 44760 10426 45152
rect 11102 44760 11162 45152
rect 11838 44760 11898 45152
rect 12574 44760 12634 45152
rect 13310 44760 13370 45152
rect 14046 44760 14106 45152
rect 14782 44760 14842 45152
rect 15518 44760 15578 45152
rect 16254 44760 16314 45152
rect 16990 44760 17050 45152
rect 17726 44760 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 640 44700 17786 44760
rect 200 9050 500 44152
rect 9800 16650 10100 44700
rect 13310 44690 13370 44700
rect 16990 44690 17050 44700
rect 9800 16649 17750 16650
rect 9800 16351 17451 16649
rect 17749 16351 17750 16649
rect 9800 16350 17750 16351
rect 200 9049 5950 9050
rect 200 8751 5651 9049
rect 5949 8751 5950 9049
rect 200 8750 5950 8751
rect 200 1000 500 8750
rect 9800 1000 10100 16350
rect 31282 1729 31462 1730
rect 31282 1551 31283 1729
rect 31461 1551 31462 1729
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 200
rect 26866 0 27046 200
rect 31282 0 31462 1551
use twin_tee_osc  twin_tee_osc_0
timestamp 1715770502
transform 1 0 138 0 1 2
box 19656 2724 30532 19940
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 4800 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 4800 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
