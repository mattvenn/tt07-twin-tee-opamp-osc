magic
tech sky130A
magscale 1 2
timestamp 1715689418
<< pwell >>
rect -201 -888 201 888
<< psubdiff >>
rect -165 818 -69 852
rect 69 818 165 852
rect -165 756 -131 818
rect 131 756 165 818
rect -165 -818 -131 -756
rect 131 -818 165 -756
rect -165 -852 -69 -818
rect 69 -852 165 -818
<< psubdiffcont >>
rect -69 818 69 852
rect -165 -756 -131 756
rect 131 -756 165 756
rect -69 -852 69 -818
<< xpolycontact >>
rect -35 290 35 722
rect -35 -722 35 -290
<< xpolyres >>
rect -35 -290 35 290
<< locali >>
rect -165 818 -69 852
rect 69 818 165 852
rect -165 756 -131 818
rect 131 756 165 818
rect -165 -818 -131 -756
rect 131 -818 165 -756
rect -165 -852 -69 -818
rect 69 -852 165 -818
<< viali >>
rect -19 307 19 704
rect -19 -704 19 -307
<< metal1 >>
rect -25 704 25 716
rect -25 307 -19 704
rect 19 307 25 704
rect -25 295 25 307
rect -25 -307 25 -295
rect -25 -704 -19 -307
rect 19 -704 25 -307
rect -25 -716 25 -704
<< properties >>
string FIXED_BBOX -148 -835 148 835
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 2.9 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 17.646k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
