** sch_path: /home/matt/work/asic-workshop/shuttle-2404/tt07-twin-tee-opamp-osc/xschem/tb_twin_tee.sch
**.subckt tb_twin_tee
V1 vdd GND 1.8
V2 vss GND 0
V3 twin_in GND 0 ac 1 0
x1 vss twin_out twin_in twin_tee
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/matt/.volare/volare/sky130/versions/bdc9412b3e468c102d01b7cf6337be06ec6e9c9a/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /home/matt/.volare/volare/sky130/versions/bdc9412b3e468c102d01b7cf6337be06ec6e9c9a/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice





.param mc_mm_switch=0
.control
ac dec 100 1 100e7
*  tran 500p 2u uic
  write testbench.raw
  set appendwrite


.endc


**** end user architecture code
**.ends

* expanding   symbol:  twin_tee.sym # of pins=3
** sym_path: /home/matt/work/asic-workshop/shuttle-2404/tt07-twin-tee-opamp-osc/xschem/twin_tee.sym
** sch_path: /home/matt/work/asic-workshop/shuttle-2404/tt07-twin-tee-opamp-osc/xschem/twin_tee.sch
.subckt twin_tee vss out in
*.iopin vss
*.iopin in
*.iopin out
XR5 c1_c2 out vss sky130_fd_pr__res_high_po_0p35 L=50 mult=1 m=1
XC1 vss c1_c2 sky130_fd_pr__cap_mim_m3_1 W=15 L=15 MF=1 m=1
XC2 vss c1_c2 sky130_fd_pr__cap_mim_m3_1 W=15 L=15 MF=1 m=1
XR4 in c1_c2 vss sky130_fd_pr__res_high_po_0p35 L=50 mult=1 m=1
XC3 in c3_c4 sky130_fd_pr__cap_mim_m3_1 W=15 L=15 MF=1 m=1
XC4 c3_c4 out sky130_fd_pr__cap_mim_m3_1 W=15 L=15 MF=1 m=1
XR6 c3_c4 vss vss sky130_fd_pr__res_high_po_0p35 L=23 mult=1 m=1
.ends

.GLOBAL GND
.end
