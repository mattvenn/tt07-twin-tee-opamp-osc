* NGSPICE file created from twin_tee_osc_parax.ext - technology: sky130A

.subckt twin_tee_osc_parax vdd vss out
X0 p3_opamp_0.VX p3_opamp_0.VBIAS.t9 vss.t36 vss.t35 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X1 vss.t7 twin_tee_0.c3_c4.t1 vss.t6 sky130_fd_pr__res_high_po_0p35 l=23
X2 vdd.t58 p3_opamp_0.V1.t7 out.t17 vdd.t57 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X3 vss.t34 p3_opamp_0.VBIAS.t10 p3_opamp_0.VX vss.t33 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X4 p3_opamp_0.VBIAS.t4 p3_opamp_0.VBIAS.t3 vss.t32 vss.t18 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=2
X5 vss.t31 p3_opamp_0.VBIAS.t5 p3_opamp_0.VBIAS.t6 vss.t18 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X6 vdd.t59 p3_opamp_0.VBIAS.t0 vss.t9 sky130_fd_pr__res_xhigh_po_0p35 l=2.9
X7 vdd.t56 p3_opamp_0.V1.t8 out.t21 vdd.t55 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X8 vdd.t2 p3_opamp_0.V2.t11 p3_opamp_0.V2.t12 vdd.t1 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=2
X9 p3_opamp_0.V2.t10 p3_opamp_0.V2.t9 vdd.t4 vdd.t3 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X10 twin_tee_0.in.t0 a_24144_17782# vss.t8 sky130_fd_pr__res_high_po_0p35 l=50.2
X11 vdd.t6 p3_opamp_0.V2.t7 p3_opamp_0.V2.t8 vdd.t5 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X12 vdd.t65 p3_opamp_0.V2.t13 p3_opamp_0.V1.t6 vdd.t64 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=2
X13 out.t19 p3_opamp_0.V1.t9 vdd.t54 vdd.t53 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X14 p3_opamp_0.VX p3_opamp_0.VBIAS.t11 vss.t30 vss.t29 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=2
X15 vdd.t0 p3_opamp_0.PLUS vss.t0 sky130_fd_pr__res_high_po_0p35 l=20
X16 vdd.t8 p3_opamp_0.V2.t14 p3_opamp_0.V1.t0 vdd.t7 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X17 p3_opamp_0.V1.t3 p3_opamp_0.V2.t15 vdd.t16 vdd.t15 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X18 vss.t26 p3_opamp_0.VBIAS.t12 p3_opamp_0.VX vss.t25 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=2
X19 out.t28 p3_opamp_0.VBIAS.t13 vss.t28 vss.t27 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=2
X20 p3_opamp_0.VBIAS.t8 p3_opamp_0.VBIAS.t7 vss.t24 vss.t18 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X21 p3_opamp_0.V2.t0 twin_tee_0.in.t1 p3_opamp_0.VX vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=0.5
X22 vdd.t52 p3_opamp_0.V1.t10 out.t15 vdd.t51 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X23 twin_tee_0.c3_c4.t2 out.t0 sky130_fd_pr__cap_mim_m3_1 l=15 w=15
X24 vdd.t50 p3_opamp_0.V1.t11 out.t8 vdd.t49 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X25 out.t27 p3_opamp_0.VBIAS.t14 vss.t23 vss.t22 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X26 vss.t21 p3_opamp_0.VBIAS.t15 out.t26 vss.t20 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X27 vss.t19 p3_opamp_0.VBIAS.t1 p3_opamp_0.VBIAS.t2 vss.t18 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=2
X28 out.t13 p3_opamp_0.V1.t12 vdd.t48 vdd.t47 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X29 vdd.t46 p3_opamp_0.V1.t13 out.t3 vdd.t45 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X30 out.t6 p3_opamp_0.V1.t14 vdd.t44 vdd.t43 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X31 vdd.t12 p3_opamp_0.V2.t5 p3_opamp_0.V2.t6 vdd.t11 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X32 vdd.t42 p3_opamp_0.V1.t15 out.t11 vdd.t41 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X33 out.t18 p3_opamp_0.V1.t16 vdd.t40 vdd.t39 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X34 p3_opamp_0.V2.t4 p3_opamp_0.V2.t3 vdd.t63 vdd.t62 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=2
X35 p3_opamp_0.V2.t2 p3_opamp_0.V2.t1 vdd.t10 vdd.t9 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X36 vdd.t38 p3_opamp_0.V1.t17 out.t4 vdd.t37 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X37 out.t12 p3_opamp_0.V1.t18 vdd.t36 vdd.t35 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X38 vdd.t14 p3_opamp_0.V2.t16 p3_opamp_0.V1.t2 vdd.t13 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X39 vdd.t34 p3_opamp_0.V1.t19 out.t20 vdd.t33 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X40 out.t5 p3_opamp_0.V1.t20 vdd.t32 vdd.t31 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X41 p3_opamp_0.V1.t4 p3_opamp_0.V2.t17 vdd.t18 vdd.t17 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X42 out.t9 p3_opamp_0.V1.t21 vdd.t30 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X43 p3_opamp_0.V1.t5 p3_opamp_0.V2.t18 vdd.t61 vdd.t60 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=2
X44 vdd.t28 p3_opamp_0.V1.t22 out.t10 vdd.t27 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X45 out.t16 p3_opamp_0.V1.t23 vdd.t26 vdd.t25 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X46 vss.t17 p3_opamp_0.VBIAS.t16 out.t25 vss.t16 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X47 out.t24 p3_opamp_0.VBIAS.t17 vss.t15 vss.t14 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X48 p3_opamp_0.V1.t1 p3_opamp_0.PLUS p3_opamp_0.VX vss.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=0.5
X49 vss.t37 a_24144_17782# sky130_fd_pr__cap_mim_m3_1 l=15 w=15
X50 out.t2 p3_opamp_0.V1.t24 vdd.t24 vdd.t23 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X51 out.t23 p3_opamp_0.VBIAS.t18 vss.t13 vss.t12 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=2
X52 vss.t11 p3_opamp_0.VBIAS.t19 out.t22 vss.t10 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X53 vss.t38 a_24144_17782# sky130_fd_pr__cap_mim_m3_1 l=15 w=15
X54 a_24144_17782# out.t1 vss.t3 sky130_fd_pr__res_high_po_0p35 l=50.2
X55 vss.t5 p3_opamp_0.PLUS vss.t4 sky130_fd_pr__res_high_po_0p35 l=20
X56 out.t7 p3_opamp_0.V1.t25 vdd.t22 vdd.t21 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X57 vdd.t20 p3_opamp_0.V1.t26 out.t14 vdd.t19 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X58 twin_tee_0.in.t2 twin_tee_0.c3_c4.t0 sky130_fd_pr__cap_mim_m3_1 l=15 w=15
R0 p3_opamp_0.VBIAS.n16 p3_opamp_0.VBIAS.n0 66.588
R1 p3_opamp_0.VBIAS.n13 p3_opamp_0.VBIAS.n1 66.588
R2 p3_opamp_0.VBIAS.n8 p3_opamp_0.VBIAS.t12 26.0899
R3 p3_opamp_0.VBIAS.n2 p3_opamp_0.VBIAS.t18 25.992
R4 p3_opamp_0.VBIAS.n7 p3_opamp_0.VBIAS.t13 25.5741
R5 p3_opamp_0.VBIAS.n11 p3_opamp_0.VBIAS.t3 25.5503
R6 p3_opamp_0.VBIAS.n14 p3_opamp_0.VBIAS.t5 25.5503
R7 p3_opamp_0.VBIAS.n15 p3_opamp_0.VBIAS.t7 25.5503
R8 p3_opamp_0.VBIAS.n17 p3_opamp_0.VBIAS.t1 25.5503
R9 p3_opamp_0.VBIAS.n2 p3_opamp_0.VBIAS.t16 25.5277
R10 p3_opamp_0.VBIAS.n3 p3_opamp_0.VBIAS.t14 25.5277
R11 p3_opamp_0.VBIAS.n4 p3_opamp_0.VBIAS.t19 25.5277
R12 p3_opamp_0.VBIAS.n5 p3_opamp_0.VBIAS.t17 25.5277
R13 p3_opamp_0.VBIAS.n6 p3_opamp_0.VBIAS.t15 25.5277
R14 p3_opamp_0.VBIAS.n8 p3_opamp_0.VBIAS.t9 25.5274
R15 p3_opamp_0.VBIAS.n9 p3_opamp_0.VBIAS.t10 25.5274
R16 p3_opamp_0.VBIAS.n10 p3_opamp_0.VBIAS.t11 25.5274
R17 p3_opamp_0.VBIAS.n0 p3_opamp_0.VBIAS.t2 17.4005
R18 p3_opamp_0.VBIAS.n0 p3_opamp_0.VBIAS.t8 17.4005
R19 p3_opamp_0.VBIAS.n1 p3_opamp_0.VBIAS.t6 17.4005
R20 p3_opamp_0.VBIAS.n1 p3_opamp_0.VBIAS.t4 17.4005
R21 p3_opamp_0.VBIAS.n12 p3_opamp_0.VBIAS.n7 7.30251
R22 p3_opamp_0.VBIAS p3_opamp_0.VBIAS.t0 3.31103
R23 p3_opamp_0.VBIAS.n11 p3_opamp_0.VBIAS.n10 1.19959
R24 p3_opamp_0.VBIAS.n10 p3_opamp_0.VBIAS.n9 0.6255
R25 p3_opamp_0.VBIAS.n9 p3_opamp_0.VBIAS.n8 0.583833
R26 p3_opamp_0.VBIAS.n3 p3_opamp_0.VBIAS.n2 0.5005
R27 p3_opamp_0.VBIAS.n5 p3_opamp_0.VBIAS.n4 0.482643
R28 p3_opamp_0.VBIAS.n6 p3_opamp_0.VBIAS.n5 0.464786
R29 p3_opamp_0.VBIAS.n4 p3_opamp_0.VBIAS.n3 0.429071
R30 p3_opamp_0.VBIAS p3_opamp_0.VBIAS.n17 0.197868
R31 p3_opamp_0.VBIAS.n15 p3_opamp_0.VBIAS.n14 0.151816
R32 p3_opamp_0.VBIAS.n7 p3_opamp_0.VBIAS.n6 0.136214
R33 p3_opamp_0.VBIAS.n14 p3_opamp_0.VBIAS.n13 0.0728684
R34 p3_opamp_0.VBIAS.n17 p3_opamp_0.VBIAS.n16 0.0728684
R35 p3_opamp_0.VBIAS.n16 p3_opamp_0.VBIAS.n15 0.0728684
R36 p3_opamp_0.VBIAS.n12 p3_opamp_0.VBIAS.n11 0.069579
R37 p3_opamp_0.VBIAS.n13 p3_opamp_0.VBIAS.n12 0.00378947
R38 vss.n64 vss.n63 258162
R39 vss.n63 vss.n62 140742
R40 vss.n65 vss.n64 92686.6
R41 vss.n63 vss.n32 21457
R42 vss.n157 vss.n151 17243.3
R43 vss.n157 vss.n152 17243.3
R44 vss.n151 vss.n6 17243.3
R45 vss.n152 vss.n6 17243.3
R46 vss.n77 vss.n43 15505.1
R47 vss.n73 vss.n43 15505.1
R48 vss.n77 vss.n44 15505.1
R49 vss.n73 vss.n44 15505.1
R50 vss.n70 vss.n46 15505.1
R51 vss.n66 vss.n46 15505.1
R52 vss.n70 vss.n47 15505.1
R53 vss.n66 vss.n47 15505.1
R54 vss.n139 vss.n7 11339.1
R55 vss.n49 vss.n7 11339.1
R56 vss.n139 vss.n8 11339.1
R57 vss.n49 vss.n8 11339.1
R58 vss.n148 vss.n141 9595.06
R59 vss.n144 vss.n141 9595.06
R60 vss.n148 vss.n142 9595.06
R61 vss.n144 vss.n142 9595.06
R62 vss.n159 vss.n2 9595.06
R63 vss.n163 vss.n2 9595.06
R64 vss.n159 vss.n3 9595.06
R65 vss.n163 vss.n3 9595.06
R66 vss.n124 vss.n29 7358.53
R67 vss.n124 vss.n30 7358.53
R68 vss.n126 vss.n30 7358.53
R69 vss.n126 vss.n29 7358.53
R70 vss.n79 vss.n35 7358.53
R71 vss.n79 vss.n36 7358.53
R72 vss.n119 vss.n36 7358.53
R73 vss.n119 vss.n35 7358.53
R74 vss.n116 vss.n38 5597.12
R75 vss.n116 vss.n39 5597.12
R76 vss.n82 vss.n38 5597.12
R77 vss.n82 vss.n39 5597.12
R78 vss.n92 vss.n89 3377.97
R79 vss.n95 vss.n89 3377.97
R80 vss.n92 vss.n90 3377.97
R81 vss.n95 vss.n90 3377.97
R82 vss.n59 vss.n51 3377.97
R83 vss.n54 vss.n51 3377.97
R84 vss.n59 vss.n52 3377.97
R85 vss.n54 vss.n52 3377.97
R86 vss.n150 vss.n140 2707.5
R87 vss.t16 vss.t12 1211.06
R88 vss.t22 vss.t16 1211.06
R89 vss.t10 vss.t22 1211.06
R90 vss.t14 vss.t10 1211.06
R91 vss.t20 vss.t14 1211.06
R92 vss.n62 vss.n50 1186.59
R93 vss.n156 vss.n153 1120.38
R94 vss.n156 vss.n155 1120.38
R95 vss.n154 vss.n153 1120.38
R96 vss.n155 vss.n154 1120.38
R97 vss.n76 vss.n45 1007.44
R98 vss.n74 vss.n45 1007.44
R99 vss.n76 vss.n75 1007.44
R100 vss.n75 vss.n74 1007.44
R101 vss.n69 vss.n48 1007.44
R102 vss.n67 vss.n48 1007.44
R103 vss.n69 vss.n68 1007.44
R104 vss.n68 vss.n67 1007.44
R105 vss.n140 vss.t12 906.971
R106 vss.t27 vss.t20 864.186
R107 vss.n80 vss.n78 855.515
R108 vss.n138 vss.n137 736.754
R109 vss.n50 vss.t27 655.605
R110 vss.n147 vss.n143 623.436
R111 vss.n145 vss.n143 623.436
R112 vss.n147 vss.n146 623.436
R113 vss.n146 vss.n145 623.436
R114 vss.n160 vss.n4 623.436
R115 vss.n162 vss.n4 623.436
R116 vss.n161 vss.n160 623.436
R117 vss.n162 vss.n161 623.436
R118 vss.n123 vss.n33 478.118
R119 vss.n137 vss.n136 451.765
R120 vss.n120 vss.n34 440.471
R121 vss.n165 vss.n164 421.781
R122 vss.n123 vss.n122 399.06
R123 vss.n138 vss.n9 399.034
R124 vss.n158 vss.t6 388.748
R125 vss.t1 vss.t33 378.079
R126 vss.n72 vss.n71 374.562
R127 vss.n152 vss.t8 373.755
R128 vss.t2 vss.t25 372.125
R129 vss.n115 vss.n40 363.671
R130 vss.n115 vss.n114 326.401
R131 vss.t2 vss.t35 309.608
R132 vss.t29 vss.t1 303.654
R133 vss.n94 vss.t29 302.166
R134 vss.t35 vss.n31 296.212
R135 vss.n68 vss.n47 292.5
R136 vss.n47 vss.t4 292.5
R137 vss.n48 vss.n46 292.5
R138 vss.n46 vss.t4 292.5
R139 vss.n75 vss.n44 292.5
R140 vss.n44 vss.t0 292.5
R141 vss.n45 vss.n43 292.5
R142 vss.n43 vss.t0 292.5
R143 vss.n114 vss.n39 292.5
R144 vss.n39 vss.t9 292.5
R145 vss.n40 vss.n38 292.5
R146 vss.n38 vss.t9 292.5
R147 vss.n155 vss.n152 292.5
R148 vss.n153 vss.n151 292.5
R149 vss.n151 vss.n150 292.5
R150 vss.n61 vss.n60 276.861
R151 vss.n60 vss.t25 233.695
R152 vss.t33 vss.n93 227.74
R153 vss.n91 vss.n87 219.482
R154 vss.n91 vss.n88 219.482
R155 vss.n96 vss.n88 219.482
R156 vss.n58 vss.n53 219.482
R157 vss.n55 vss.n53 219.482
R158 vss.n56 vss.n55 219.482
R159 vss.n118 vss.n37 215.702
R160 vss.n122 vss.n120 208.189
R161 vss.n55 vss.n54 195
R162 vss.n54 vss.n31 195
R163 vss.n59 vss.n58 195
R164 vss.n60 vss.n59 195
R165 vss.n96 vss.n95 195
R166 vss.n95 vss.n94 195
R167 vss.n92 vss.n91 195
R168 vss.n93 vss.n92 195
R169 vss.n94 vss.n37 165.083
R170 vss.t6 vss.n5 159.375
R171 vss.n57 vss.n56 134.776
R172 vss.n18 vss.n9 130.133
R173 vss.n97 vss.n87 128
R174 vss.n35 vss.n34 117.001
R175 vss.t18 vss.n35 117.001
R176 vss.n49 vss.n10 117.001
R177 vss.n50 vss.n49 117.001
R178 vss.n139 vss.n138 117.001
R179 vss.n140 vss.n139 117.001
R180 vss.n33 vss.n29 117.001
R181 vss.n61 vss.n29 117.001
R182 vss.n121 vss.n30 117.001
R183 vss.n37 vss.n30 117.001
R184 vss.n102 vss.n36 117.001
R185 vss.t18 vss.n36 117.001
R186 vss.n27 vss.n11 110.359
R187 vss.n117 vss.t9 107.85
R188 vss.n78 vss.t0 107.85
R189 vss.n72 vss.t0 107.85
R190 vss.n71 vss.t4 107.85
R191 vss.n65 vss.t4 107.85
R192 vss.n81 vss.t18 107.123
R193 vss.n97 vss.n96 91.4829
R194 vss.n109 vss.t32 86.2761
R195 vss.n108 vss.t19 86.2684
R196 vss.n16 vss.t28 86.2495
R197 vss.n23 vss.t26 85.2172
R198 vss.n98 vss.t30 85.2172
R199 vss.n93 vss.n32 84.8449
R200 vss.n84 vss.n40 81.1864
R201 vss.n81 vss.n80 80.1595
R202 vss.n118 vss.n117 78.7021
R203 vss.n58 vss.n57 78.0993
R204 vss.n21 vss.n11 73.4123
R205 vss.n130 vss.n24 68.9308
R206 vss.n14 vss.n13 68.8514
R207 vss.n62 vss.n61 68.4714
R208 vss.n108 vss.n107 68.1549
R209 vss.n16 vss.n15 68.0911
R210 vss.n14 vss.n12 68.0905
R211 vss.n64 vss.t8 65.8985
R212 vss.n149 vss.t3 58.5301
R213 vss.t3 vss.n5 58.5301
R214 vss.n158 vss.t8 58.5301
R215 vss.n164 vss.t8 58.5301
R216 vss.n56 vss.n52 58.5005
R217 vss.n52 vss.t2 58.5005
R218 vss.n53 vss.n51 58.5005
R219 vss.t2 vss.n51 58.5005
R220 vss.n90 vss.n87 58.5005
R221 vss.t1 vss.n90 58.5005
R222 vss.n89 vss.n88 58.5005
R223 vss.t1 vss.n89 58.5005
R224 vss.n102 vss.n42 55.9122
R225 vss.n163 vss.n162 48.7505
R226 vss.n164 vss.n163 48.7505
R227 vss.n160 vss.n159 48.7505
R228 vss.n159 vss.n158 48.7505
R229 vss.n145 vss.n144 48.7505
R230 vss.n144 vss.n5 48.7505
R231 vss.n148 vss.n147 48.7505
R232 vss.n149 vss.n148 48.7505
R233 vss.n113 vss.n112 45.5155
R234 vss.n125 vss.n31 44.6554
R235 vss.n104 vss.t7 44.1758
R236 vss.n105 vss.t5 43.3392
R237 vss.n127 vss.n28 33.5081
R238 vss.n113 vss.n41 30.6245
R239 vss.n125 vss.n32 28.282
R240 vss.n116 vss.n115 26.5914
R241 vss.n117 vss.n116 26.5914
R242 vss.n83 vss.n82 26.5914
R243 vss.n82 vss.n81 26.5914
R244 vss.n18 vss.n10 23.8938
R245 vss.n150 vss.n149 22.1468
R246 vss.n124 vss.n123 20.8934
R247 vss.n125 vss.n124 20.8934
R248 vss.n120 vss.n119 20.8934
R249 vss.n119 vss.n118 20.8934
R250 vss.n127 vss.n126 20.8934
R251 vss.n126 vss.n125 20.8934
R252 vss.n79 vss.n42 20.8934
R253 vss.n80 vss.n79 20.8934
R254 vss.n161 vss.n3 17.7278
R255 vss.n3 vss.t8 17.7278
R256 vss.n4 vss.n2 17.7278
R257 vss.n2 vss.t8 17.7278
R258 vss.n146 vss.n142 17.7278
R259 vss.n142 vss.t3 17.7278
R260 vss.n143 vss.n141 17.7278
R261 vss.n141 vss.t3 17.7278
R262 vss.n107 vss.t24 17.4005
R263 vss.n107 vss.t31 17.4005
R264 vss.n24 vss.t36 17.4005
R265 vss.n24 vss.t34 17.4005
R266 vss.n15 vss.t15 17.4005
R267 vss.n15 vss.t21 17.4005
R268 vss.n12 vss.t23 17.4005
R269 vss.n12 vss.t11 17.4005
R270 vss.n13 vss.t13 17.4005
R271 vss.n13 vss.t17 17.4005
R272 vss.n135 vss.n11 13.6763
R273 vss.n128 vss.n27 12.5161
R274 vss.n9 vss.n7 12.188
R275 vss.t10 vss.n7 12.188
R276 vss.n137 vss.n8 12.188
R277 vss.t10 vss.n8 12.188
R278 vss.n102 vss.n28 11.6757
R279 vss.n84 vss.n83 9.6645
R280 vss.n121 vss.n28 9.30959
R281 vss.n122 vss.n121 8.14595
R282 vss.n67 vss.n66 8.0142
R283 vss.n66 vss.n65 8.0142
R284 vss.n70 vss.n69 8.0142
R285 vss.n71 vss.n70 8.0142
R286 vss.n74 vss.n73 8.0142
R287 vss.n73 vss.n72 8.0142
R288 vss.n77 vss.n76 8.0142
R289 vss.n78 vss.n77 8.0142
R290 vss.n33 vss.n21 7.52991
R291 vss.n114 vss.n113 7.51354
R292 vss.n113 vss.n34 7.51354
R293 vss.n154 vss.n6 7.22272
R294 vss.t6 vss.n6 7.22272
R295 vss.n157 vss.n156 7.22272
R296 vss.t6 vss.n157 7.22272
R297 vss.n136 vss.n10 7.05622
R298 vss.n98 vss.n97 6.55702
R299 vss.n57 vss.n23 6.54313
R300 vss.n101 vss.n100 4.50397
R301 vss.n132 vss.n131 4.5005
R302 vss.n130 vss.n129 4.5005
R303 vss.n112 vss.n42 4.06119
R304 vss.n106 vss.n105 4.00099
R305 vss.n135 vss.n134 3.16116
R306 vss.n19 vss.n18 3.1005
R307 vss.n133 vss.n21 2.42272
R308 vss.n1 vss.n0 2.10264
R309 vss.n104 vss.n1 2.04087
R310 vss.n103 vss.n102 1.8605
R311 vss.n20 vss.n10 1.5505
R312 vss.n19 vss.n17 1.30682
R313 vss.n165 vss.n1 1.27326
R314 vss.n105 vss.n104 0.943777
R315 vss.n0 vss.t38 0.894893
R316 vss.t18 vss.t9 0.729218
R317 vss.n111 vss.n85 0.69889
R318 vss.n100 vss.n99 0.628972
R319 vss.n131 vss.n130 0.622028
R320 vss.n85 vss.n84 0.554989
R321 vss.n17 vss.n16 0.504667
R322 vss.n85 vss.n41 0.4655
R323 vss.n166 vss 0.441333
R324 vss.n83 vss.n41 0.4165
R325 vss.n110 vss.n106 0.379288
R326 vss.n112 vss.n111 0.358192
R327 vss.n129 vss.n128 0.344944
R328 vss.n131 vss.n23 0.311665
R329 vss.n100 vss.n98 0.308192
R330 vss vss.n166 0.274878
R331 vss.n17 vss.n14 0.263
R332 vss.n101 vss.n86 0.242521
R333 vss.n134 vss.n133 0.211936
R334 vss.n20 vss.n19 0.202941
R335 vss.n103 vss.n101 0.170929
R336 vss.n99 vss.n86 0.1505
R337 vss.n26 vss.n25 0.1505
R338 vss.n132 vss.n22 0.121511
R339 vss.n129 vss.n22 0.117521
R340 vss.n136 vss.n135 0.108289
R341 vss.n134 vss.n20 0.106883
R342 vss.n0 vss.t37 0.0927731
R343 vss.n27 vss.n22 0.0882358
R344 vss vss.n103 0.0866169
R345 vss.n110 vss.n109 0.0755
R346 vss.n133 vss.n132 0.063
R347 vss.n128 vss.n127 0.0573889
R348 vss vss.n165 0.0479585
R349 vss.n111 vss.n110 0.032697
R350 vss.n130 vss.n25 0.0143889
R351 vss.n106 vss 0.013548
R352 vss.n166 vss 0.0119108
R353 vss.n129 vss.n26 0.00581915
R354 vss.n109 vss.n108 0.00440625
R355 vss.n99 vss.n25 0.00397222
R356 vss.n86 vss.n26 0.00182979
R357 twin_tee_0.c3_c4 twin_tee_0.c3_c4.t1 46.7014
R358 twin_tee_0.c3_c4 twin_tee_0.c3_c4.t0 0.349462
R359 twin_tee_0.c3_c4 twin_tee_0.c3_c4.n0 0.0354413
R360 twin_tee_0.c3_c4.n0 twin_tee_0.c3_c4.t2 0.0274722
R361 twin_tee_0.c3_c4.n0 twin_tee_0.c3_c4 0.0109069
R362 p3_opamp_0.V1.n1 p3_opamp_0.V1.t8 240.631
R363 p3_opamp_0.V1.n0 p3_opamp_0.V1.t20 240.631
R364 p3_opamp_0.V1.n0 p3_opamp_0.V1.t7 240.349
R365 p3_opamp_0.V1.n0 p3_opamp_0.V1.t24 240.349
R366 p3_opamp_0.V1.n1 p3_opamp_0.V1.t16 240.349
R367 p3_opamp_0.V1.n1 p3_opamp_0.V1.t10 240.349
R368 p3_opamp_0.V1.n1 p3_opamp_0.V1.t12 240.349
R369 p3_opamp_0.V1.n1 p3_opamp_0.V1.t13 240.349
R370 p3_opamp_0.V1.n1 p3_opamp_0.V1.t9 240.349
R371 p3_opamp_0.V1.n1 p3_opamp_0.V1.t22 240.349
R372 p3_opamp_0.V1.n1 p3_opamp_0.V1.t14 240.349
R373 p3_opamp_0.V1.n0 p3_opamp_0.V1.t17 240.349
R374 p3_opamp_0.V1.n0 p3_opamp_0.V1.t21 240.349
R375 p3_opamp_0.V1.n0 p3_opamp_0.V1.t11 240.349
R376 p3_opamp_0.V1.n0 p3_opamp_0.V1.t25 240.349
R377 p3_opamp_0.V1.n0 p3_opamp_0.V1.t19 240.349
R378 p3_opamp_0.V1.n0 p3_opamp_0.V1.t23 240.349
R379 p3_opamp_0.V1.n0 p3_opamp_0.V1.t15 240.349
R380 p3_opamp_0.V1.n0 p3_opamp_0.V1.t18 240.349
R381 p3_opamp_0.V1.n0 p3_opamp_0.V1.t26 240.349
R382 p3_opamp_0.V1 p3_opamp_0.V1.t5 230.536
R383 p3_opamp_0.V1.n4 p3_opamp_0.V1.t6 229.337
R384 p3_opamp_0.V1 p3_opamp_0.V1.n3 201.905
R385 p3_opamp_0.V1 p3_opamp_0.V1.n2 201.904
R386 p3_opamp_0.V1.n4 p3_opamp_0.V1.t1 36.1494
R387 p3_opamp_0.V1.n3 p3_opamp_0.V1.t0 28.5655
R388 p3_opamp_0.V1.n3 p3_opamp_0.V1.t4 28.5655
R389 p3_opamp_0.V1.n2 p3_opamp_0.V1.t2 28.5655
R390 p3_opamp_0.V1.n2 p3_opamp_0.V1.t3 28.5655
R391 p3_opamp_0.V1 p3_opamp_0.V1.n0 8.1351
R392 p3_opamp_0.V1 p3_opamp_0.V1.n4 4.80549
R393 p3_opamp_0.V1.n0 p3_opamp_0.V1.n1 4.75675
R394 out.n6 out.n5 203.756
R395 out.n6 out.n4 203.499
R396 out.n28 out.n8 201.875
R397 out.n27 out.n9 201.695
R398 out.n24 out.n12 201.619
R399 out.n22 out.n14 201.619
R400 out.n23 out.n13 201.619
R401 out.n26 out.n10 201.619
R402 out.n19 out.n17 201.561
R403 out.n20 out.n16 201.561
R404 out.n7 out.t23 83.7297
R405 out.n19 out.n18 69.1449
R406 out.n21 out.n15 68.1265
R407 out.n25 out.n11 68.1259
R408 out.n0 out.t1 44.2614
R409 out.n12 out.t8 28.5655
R410 out.n12 out.t7 28.5655
R411 out.n17 out.t14 28.5655
R412 out.n17 out.t5 28.5655
R413 out.n16 out.t17 28.5655
R414 out.n16 out.t2 28.5655
R415 out.n14 out.t11 28.5655
R416 out.n14 out.t12 28.5655
R417 out.n13 out.t20 28.5655
R418 out.n13 out.t16 28.5655
R419 out.n10 out.t4 28.5655
R420 out.n10 out.t9 28.5655
R421 out.n9 out.t10 28.5655
R422 out.n9 out.t6 28.5655
R423 out.n8 out.t3 28.5655
R424 out.n8 out.t19 28.5655
R425 out.n5 out.t15 28.5655
R426 out.n5 out.t13 28.5655
R427 out.n4 out.t21 28.5655
R428 out.n4 out.t18 28.5655
R429 out.n11 out.t25 17.4005
R430 out.n11 out.t27 17.4005
R431 out.n15 out.t22 17.4005
R432 out.n15 out.t24 17.4005
R433 out.n18 out.t26 17.4005
R434 out.n18 out.t28 17.4005
R435 out.n0 out.t0 4.93405
R436 out.n31 out.n2 2.69072
R437 out.n2 out 2.15883
R438 out.n29 out.n7 1.38826
R439 out.n30 out.n29 0.663586
R440 out.n24 out 0.565168
R441 out.n29 out.n28 0.285222
R442 out.n2 out.n1 0.17767
R443 out.n23 out.n22 0.154346
R444 out.n27 out.n26 0.151942
R445 out.n24 out.n23 0.149538
R446 out.n20 out.n19 0.149538
R447 out.n26 out.n25 0.139923
R448 out.n28 out.n27 0.1255
R449 out.n22 out.n21 0.1255
R450 out out.n31 0.1255
R451 out out.n30 0.0929762
R452 out.n1 out 0.0713874
R453 out.n29 out.n6 0.0639766
R454 out.n30 out.n3 0.0635409
R455 out.n31 out 0.063
R456 out.n1 out 0.0609244
R457 out.n21 out.n20 0.0269423
R458 out out.n3 0.0264615
R459 out out.n0 0.0167338
R460 out.n25 out.n24 0.0149231
R461 out.n7 out.n3 0.00499257
R462 vdd.n50 vdd.n45 6857.65
R463 vdd.n50 vdd.n46 6857.65
R464 vdd.n48 vdd.n46 6857.65
R465 vdd.n48 vdd.n45 6857.65
R466 vdd.n11 vdd.n6 6130.59
R467 vdd.n11 vdd.n7 6130.59
R468 vdd.n9 vdd.n7 6130.59
R469 vdd.n9 vdd.n6 6130.59
R470 vdd.n25 vdd.n22 6130.59
R471 vdd.n25 vdd.n23 6130.59
R472 vdd.n27 vdd.n23 6130.59
R473 vdd.n27 vdd.n22 6130.59
R474 vdd.n47 vdd.n43 731.482
R475 vdd.n47 vdd.n44 731.482
R476 vdd.t5 vdd.t62 681.976
R477 vdd.t9 vdd.t5 681.976
R478 vdd.t11 vdd.t3 681.976
R479 vdd.t3 vdd.t1 681.976
R480 vdd.t7 vdd.t60 681.976
R481 vdd.t17 vdd.t7 681.976
R482 vdd.t13 vdd.t15 681.976
R483 vdd.t15 vdd.t64 681.976
R484 vdd.n8 vdd.n4 653.929
R485 vdd.n8 vdd.n5 653.929
R486 vdd.n24 vdd.n20 653.929
R487 vdd.n24 vdd.n21 653.929
R488 vdd.n51 vdd.n44 646.381
R489 vdd.n52 vdd.n43 625.601
R490 vdd.t62 vdd.n6 541.571
R491 vdd.t1 vdd.n7 541.571
R492 vdd.t60 vdd.n22 541.571
R493 vdd.t64 vdd.n23 541.571
R494 vdd.n12 vdd.n5 493.892
R495 vdd.n28 vdd.n21 487.142
R496 vdd.n13 vdd.n4 381.115
R497 vdd.n29 vdd.n20 372.925
R498 vdd.n10 vdd.t9 340.988
R499 vdd.n10 vdd.t11 340.988
R500 vdd.n26 vdd.t17 340.988
R501 vdd.n26 vdd.t13 340.988
R502 vdd.t55 vdd.n45 318.216
R503 vdd.t31 vdd.n46 318.216
R504 vdd.t39 vdd.t55 235.267
R505 vdd.t51 vdd.t39 235.267
R506 vdd.t47 vdd.t51 235.267
R507 vdd.t45 vdd.t47 235.267
R508 vdd.t53 vdd.t45 235.267
R509 vdd.t27 vdd.t53 235.267
R510 vdd.t43 vdd.t27 235.267
R511 vdd.t37 vdd.t43 235.267
R512 vdd.t29 vdd.t37 235.267
R513 vdd.t49 vdd.t21 235.267
R514 vdd.t21 vdd.t33 235.267
R515 vdd.t33 vdd.t25 235.267
R516 vdd.t25 vdd.t41 235.267
R517 vdd.t41 vdd.t35 235.267
R518 vdd.t35 vdd.t57 235.267
R519 vdd.t57 vdd.t23 235.267
R520 vdd.t23 vdd.t19 235.267
R521 vdd.t19 vdd.t31 235.267
R522 vdd.n34 vdd.t56 230.56
R523 vdd.n60 vdd.t32 230.405
R524 vdd.n15 vdd.n3 202.125
R525 vdd.n18 vdd.n1 201.834
R526 vdd.n16 vdd.n2 201.834
R527 vdd.n65 vdd.n56 201.779
R528 vdd.n35 vdd.n32 201.779
R529 vdd.n70 vdd.n41 201.761
R530 vdd.n34 vdd.n33 201.761
R531 vdd.n74 vdd.n37 201.761
R532 vdd.n73 vdd.n38 201.761
R533 vdd.n71 vdd.n40 201.761
R534 vdd.n66 vdd.n55 201.756
R535 vdd.n36 vdd.n31 201.756
R536 vdd.n63 vdd.n57 201.744
R537 vdd.n59 vdd.n58 201.744
R538 vdd.n72 vdd.n39 201.704
R539 vdd.n49 vdd.t29 117.633
R540 vdd.n49 vdd.t49 117.633
R541 vdd.n13 vdd.n12 44.5872
R542 vdd.n29 vdd.n28 43.1489
R543 vdd.n79 vdd.t0 43.0539
R544 vdd.n78 vdd.t59 42.7092
R545 vdd.n6 vdd.n4 30.8338
R546 vdd.n7 vdd.n5 30.8338
R547 vdd.n22 vdd.n20 30.8338
R548 vdd.n23 vdd.n21 30.8338
R549 vdd.n45 vdd.n43 30.8338
R550 vdd.n46 vdd.n44 30.8338
R551 vdd.n1 vdd.t63 28.5655
R552 vdd.n1 vdd.t6 28.5655
R553 vdd.n2 vdd.t10 28.5655
R554 vdd.n2 vdd.t12 28.5655
R555 vdd.n3 vdd.t4 28.5655
R556 vdd.n3 vdd.t2 28.5655
R557 vdd.n41 vdd.t22 28.5655
R558 vdd.n41 vdd.t34 28.5655
R559 vdd.n55 vdd.t26 28.5655
R560 vdd.n55 vdd.t42 28.5655
R561 vdd.n57 vdd.t36 28.5655
R562 vdd.n57 vdd.t58 28.5655
R563 vdd.n58 vdd.t24 28.5655
R564 vdd.n58 vdd.t20 28.5655
R565 vdd.n56 vdd.t16 28.5655
R566 vdd.n56 vdd.t65 28.5655
R567 vdd.n39 vdd.t18 28.5655
R568 vdd.n39 vdd.t14 28.5655
R569 vdd.n32 vdd.t61 28.5655
R570 vdd.n32 vdd.t8 28.5655
R571 vdd.n33 vdd.t40 28.5655
R572 vdd.n33 vdd.t52 28.5655
R573 vdd.n31 vdd.t48 28.5655
R574 vdd.n31 vdd.t46 28.5655
R575 vdd.n37 vdd.t54 28.5655
R576 vdd.n37 vdd.t28 28.5655
R577 vdd.n38 vdd.t44 28.5655
R578 vdd.n38 vdd.t38 28.5655
R579 vdd.n40 vdd.t30 28.5655
R580 vdd.n40 vdd.t50 28.5655
R581 vdd.n52 vdd.n51 15.3605
R582 vdd.n9 vdd.n8 4.5127
R583 vdd.n10 vdd.n9 4.5127
R584 vdd.n12 vdd.n11 4.5127
R585 vdd.n11 vdd.n10 4.5127
R586 vdd.n25 vdd.n24 4.5127
R587 vdd.n26 vdd.n25 4.5127
R588 vdd.n28 vdd.n27 4.5127
R589 vdd.n27 vdd.n26 4.5127
R590 vdd.n48 vdd.n47 3.85467
R591 vdd.n49 vdd.n48 3.85467
R592 vdd.n51 vdd.n50 3.85467
R593 vdd.n50 vdd.n49 3.85467
R594 vdd.n79 vdd 2.02508
R595 vdd.n67 vdd.n66 1.5005
R596 vdd.n70 vdd.n69 1.5005
R597 vdd.n61 vdd.n60 1.01532
R598 vdd.n19 vdd.n18 0.903037
R599 vdd.n77 vdd.n76 0.82517
R600 vdd.n68 vdd.n42 0.7505
R601 vdd.n64 vdd.n54 0.7505
R602 vdd vdd.n79 0.521599
R603 vdd.n18 vdd.n17 0.338735
R604 vdd.n17 vdd.n16 0.338735
R605 vdd.n14 vdd.n13 0.282318
R606 vdd.n30 vdd.n29 0.282318
R607 vdd.n15 vdd.n14 0.275967
R608 vdd.n16 vdd.n15 0.256696
R609 vdd.n74 vdd.n73 0.235794
R610 vdd.n71 vdd.n70 0.235794
R611 vdd.n53 vdd.n52 0.216779
R612 vdd.n75 vdd.n36 0.195353
R613 vdd.n77 vdd.n19 0.195317
R614 vdd.n60 vdd.n59 0.191472
R615 vdd.n63 vdd.n62 0.181056
R616 vdd.n19 vdd.n0 0.174399
R617 vdd.n17 vdd.n0 0.173577
R618 vdd.n62 vdd.n61 0.167167
R619 vdd.n61 vdd.n54 0.137765
R620 vdd.n35 vdd.n34 0.136529
R621 vdd.n78 vdd.n77 0.136138
R622 vdd.n72 vdd.n71 0.118147
R623 vdd.n64 vdd.n63 0.116513
R624 vdd.n70 vdd.n42 0.114471
R625 vdd.n66 vdd.n42 0.114471
R626 vdd.n73 vdd.n72 0.110794
R627 vdd.n69 vdd.n53 0.0996848
R628 vdd.n36 vdd.n35 0.0924118
R629 vdd.n66 vdd.n65 0.0924118
R630 vdd.n14 vdd.n0 0.0897857
R631 vdd.n76 vdd.n30 0.0888152
R632 vdd.n53 vdd.n30 0.0860978
R633 vdd.n76 vdd.n75 0.0755
R634 vdd vdd.n78 0.063
R635 vdd.n67 vdd.n54 0.0439783
R636 vdd.n69 vdd.n68 0.0426196
R637 vdd.n68 vdd.n67 0.0426196
R638 vdd.n62 vdd.n59 0.0421667
R639 vdd.n75 vdd.n74 0.0409412
R640 vdd.n65 vdd.n64 0.0262353
R641 p3_opamp_0.V2 p3_opamp_0.V2.t12 228.542
R642 p3_opamp_0.V2 p3_opamp_0.V2.t4 228.456
R643 p3_opamp_0.V2 p3_opamp_0.V2.n0 199.977
R644 p3_opamp_0.V2 p3_opamp_0.V2.n1 199.923
R645 p3_opamp_0.V2 p3_opamp_0.V2.t0 34.7182
R646 p3_opamp_0.V2.n0 p3_opamp_0.V2.t6 28.5655
R647 p3_opamp_0.V2.n0 p3_opamp_0.V2.t10 28.5655
R648 p3_opamp_0.V2.n1 p3_opamp_0.V2.t8 28.5655
R649 p3_opamp_0.V2.n1 p3_opamp_0.V2.t2 28.5655
R650 p3_opamp_0.V2 p3_opamp_0.V2.t3 26.6205
R651 p3_opamp_0.V2 p3_opamp_0.V2.t18 26.0942
R652 p3_opamp_0.V2 p3_opamp_0.V2.t14 26.0942
R653 p3_opamp_0.V2 p3_opamp_0.V2.t17 26.0942
R654 p3_opamp_0.V2 p3_opamp_0.V2.t16 26.0942
R655 p3_opamp_0.V2 p3_opamp_0.V2.t15 26.0942
R656 p3_opamp_0.V2 p3_opamp_0.V2.t13 26.0942
R657 p3_opamp_0.V2 p3_opamp_0.V2.t11 26.05
R658 p3_opamp_0.V2 p3_opamp_0.V2.t9 26.05
R659 p3_opamp_0.V2 p3_opamp_0.V2.t5 26.0489
R660 p3_opamp_0.V2 p3_opamp_0.V2.t1 26.0488
R661 p3_opamp_0.V2 p3_opamp_0.V2.t7 26.0478
R662 twin_tee_0.in.n2 twin_tee_0.in.t1 154.407
R663 twin_tee_0.in.n0 twin_tee_0.in.t0 43.1124
R664 twin_tee_0.in.n0 twin_tee_0.in.t2 10.2463
R665 twin_tee_0.in twin_tee_0.in.n5 9.43796
R666 twin_tee_0.in.n5 twin_tee_0.in.n4 4.5005
R667 twin_tee_0.in.n3 twin_tee_0.in.n1 2.2505
R668 twin_tee_0.in.n2 twin_tee_0.in.n1 1.48465
R669 twin_tee_0.in twin_tee_0.in.n0 0.723459
R670 twin_tee_0.in.n4 twin_tee_0.in.n2 0.394718
R671 twin_tee_0.in.n3 twin_tee_0.in 0.054875
R672 twin_tee_0.in.n5 twin_tee_0.in.n1 0.0307083
R673 twin_tee_0.in.n4 twin_tee_0.in.n3 0.002375
C0 p3_opamp_0.V2 p3_opamp_0.VBIAS 0.190761f
C1 out twin_tee_0.c3_c4 21.970499f
C2 p3_opamp_0.V2 out 0.004966f
C3 p3_opamp_0.V1 vdd 9.40784f
C4 p3_opamp_0.VX twin_tee_0.in 0.578867f
C5 p3_opamp_0.V1 twin_tee_0.in 0.01158f
C6 out p3_opamp_0.VBIAS 2.97334f
C7 vdd twin_tee_0.c3_c4 0.280465f
C8 p3_opamp_0.V2 vdd 14.0343f
C9 twin_tee_0.in twin_tee_0.c3_c4 21.3079f
C10 p3_opamp_0.VX p3_opamp_0.PLUS 0.579422f
C11 p3_opamp_0.V1 p3_opamp_0.PLUS 0.654269f
C12 p3_opamp_0.V2 twin_tee_0.in 0.55445f
C13 vdd p3_opamp_0.VBIAS 0.904071f
C14 twin_tee_0.in p3_opamp_0.VBIAS 0.71001f
C15 out vdd 5.12667f
C16 p3_opamp_0.V2 p3_opamp_0.PLUS 0.04754f
C17 a_24144_17782# twin_tee_0.c3_c4 0.257745f
C18 p3_opamp_0.PLUS p3_opamp_0.VBIAS 0.738369f
C19 out p3_opamp_0.PLUS 0.455883f
C20 vdd twin_tee_0.in 0.53616f
C21 out a_24144_17782# 1.17749f
C22 vdd p3_opamp_0.PLUS 0.52756f
C23 p3_opamp_0.V1 p3_opamp_0.VX 0.096512f
C24 twin_tee_0.in p3_opamp_0.PLUS 0.041f
C25 a_24144_17782# twin_tee_0.in 1.64671f
C26 p3_opamp_0.V1 twin_tee_0.c3_c4 0.011866f
C27 p3_opamp_0.V2 p3_opamp_0.VX 0.119464f
C28 p3_opamp_0.V2 p3_opamp_0.V1 6.83344f
C29 p3_opamp_0.VX p3_opamp_0.VBIAS 1.88665f
C30 p3_opamp_0.V1 p3_opamp_0.VBIAS 0.241132f
C31 p3_opamp_0.V2 twin_tee_0.c3_c4 0.010504f
C32 out p3_opamp_0.VX 1.32e-21
C33 p3_opamp_0.V1 out 2.01513f
C34 out vss 16.742512f
C35 vdd vss 34.76403f
C36 p3_opamp_0.VX vss 1.45094f
C37 p3_opamp_0.V1 vss 12.799731f
C38 p3_opamp_0.V2 vss 21.569592f
C39 p3_opamp_0.VBIAS vss 26.706236f
C40 p3_opamp_0.PLUS vss 8.79069f
C41 twin_tee_0.c3_c4 vss 9.77696f
C42 twin_tee_0.in vss 21.124464f
C43 a_24144_17782# vss 57.9734f
C44 twin_tee_0.in.t2 vss 16.2946f
C45 twin_tee_0.in.t0 vss 0.010986f
C46 twin_tee_0.in.n0 vss 0.979236f
C47 twin_tee_0.in.n1 vss 0.097937f
C48 twin_tee_0.in.t1 vss 0.045094f
C49 twin_tee_0.in.n2 vss 0.0445f
C50 twin_tee_0.in.n3 vss 0.008073f
C51 twin_tee_0.in.n4 vss 0.033356f
C52 twin_tee_0.in.n5 vss 1.40238f
C53 p3_opamp_0.V2.t0 vss 0.093093f
C54 p3_opamp_0.V2.t13 vss 0.456467f
C55 p3_opamp_0.V2.t12 vss 0.039293f
C56 p3_opamp_0.V2.t6 vss 0.01067f
C57 p3_opamp_0.V2.t10 vss 0.01067f
C58 p3_opamp_0.V2.n0 vss 0.022041f
C59 p3_opamp_0.V2.t8 vss 0.01067f
C60 p3_opamp_0.V2.t2 vss 0.01067f
C61 p3_opamp_0.V2.n1 vss 0.022034f
C62 p3_opamp_0.V2.t18 vss 0.456467f
C63 p3_opamp_0.V2.t14 vss 0.456467f
C64 p3_opamp_0.V2.t17 vss 0.456467f
C65 p3_opamp_0.V2.t16 vss 0.456467f
C66 p3_opamp_0.V2.t15 vss 0.456467f
C67 p3_opamp_0.V2.t4 vss 0.039293f
C68 p3_opamp_0.V2.t3 vss 0.45557f
C69 p3_opamp_0.V2.t7 vss 0.455564f
C70 p3_opamp_0.V2.t1 vss 0.45557f
C71 p3_opamp_0.V2.t5 vss 0.45557f
C72 p3_opamp_0.V2.t9 vss 0.45557f
C73 p3_opamp_0.V2.t11 vss 0.45557f
C74 vdd.t59 vss 0.019809f
C75 vdd.n0 vss 0.223596f
C76 vdd.t63 vss 0.005014f
C77 vdd.t6 vss 0.005014f
C78 vdd.n1 vss 0.010764f
C79 vdd.t10 vss 0.005014f
C80 vdd.t12 vss 0.005014f
C81 vdd.n2 vss 0.010764f
C82 vdd.t4 vss 0.005014f
C83 vdd.t2 vss 0.005014f
C84 vdd.n3 vss 0.011133f
C85 vdd.n4 vss 0.110301f
C86 vdd.n5 vss 0.105891f
C87 vdd.n6 vss 0.337331f
C88 vdd.n7 vss 0.337331f
C89 vdd.t62 vss 0.455865f
C90 vdd.t5 vss 0.505191f
C91 vdd.t9 vss 0.378893f
C92 vdd.t1 vss 0.455865f
C93 vdd.t3 vss 0.505191f
C94 vdd.t11 vss 0.378893f
C95 vdd.n8 vss 0.102411f
C96 vdd.n9 vss 0.102411f
C97 vdd.n10 vss 0.252596f
C98 vdd.n11 vss 0.102411f
C99 vdd.n12 vss 0.10405f
C100 vdd.n13 vss 0.096749f
C101 vdd.n14 vss 0.427321f
C102 vdd.n15 vss 0.676018f
C103 vdd.n16 vss 0.22694f
C104 vdd.n17 vss 0.1352f
C105 vdd.n18 vss 0.180024f
C106 vdd.n19 vss 0.310158f
C107 vdd.n20 vss 0.111125f
C108 vdd.n21 vss 0.10601f
C109 vdd.n22 vss 0.337331f
C110 vdd.n23 vss 0.337331f
C111 vdd.t60 vss 0.455865f
C112 vdd.t7 vss 0.505191f
C113 vdd.t17 vss 0.378893f
C114 vdd.n24 vss 0.102411f
C115 vdd.n25 vss 0.102411f
C116 vdd.t64 vss 0.455865f
C117 vdd.t15 vss 0.505191f
C118 vdd.t13 vss 0.378893f
C119 vdd.n26 vss 0.252596f
C120 vdd.n27 vss 0.102411f
C121 vdd.n28 vss 0.107685f
C122 vdd.n29 vss 0.100401f
C123 vdd.n30 vss 0.254494f
C124 vdd.t48 vss 0.005014f
C125 vdd.t46 vss 0.005014f
C126 vdd.n31 vss 0.010787f
C127 vdd.t61 vss 0.005014f
C128 vdd.t8 vss 0.005014f
C129 vdd.n32 vss 0.010772f
C130 vdd.t40 vss 0.005014f
C131 vdd.t52 vss 0.005014f
C132 vdd.n33 vss 0.010787f
C133 vdd.t56 vss 0.019032f
C134 vdd.n34 vss 0.348583f
C135 vdd.n35 vss 0.135105f
C136 vdd.n36 vss 0.158338f
C137 vdd.t54 vss 0.005014f
C138 vdd.t28 vss 0.005014f
C139 vdd.n37 vss 0.010787f
C140 vdd.t44 vss 0.005014f
C141 vdd.t38 vss 0.005014f
C142 vdd.n38 vss 0.010783f
C143 vdd.t18 vss 0.005014f
C144 vdd.t14 vss 0.005014f
C145 vdd.n39 vss 0.010759f
C146 vdd.t30 vss 0.005014f
C147 vdd.t50 vss 0.005014f
C148 vdd.n40 vss 0.010783f
C149 vdd.t22 vss 0.005014f
C150 vdd.t34 vss 0.005014f
C151 vdd.n41 vss 0.010787f
C152 vdd.n42 vss 0.045557f
C153 vdd.n43 vss 0.119518f
C154 vdd.n44 vss 0.120066f
C155 vdd.n45 vss 0.264865f
C156 vdd.n46 vss 0.264865f
C157 vdd.t55 vss 0.209561f
C158 vdd.t39 vss 0.17428f
C159 vdd.t51 vss 0.17428f
C160 vdd.t47 vss 0.17428f
C161 vdd.t45 vss 0.17428f
C162 vdd.t53 vss 0.17428f
C163 vdd.t27 vss 0.17428f
C164 vdd.t43 vss 0.17428f
C165 vdd.t37 vss 0.17428f
C166 vdd.t29 vss 0.13071f
C167 vdd.t31 vss 0.209561f
C168 vdd.t19 vss 0.17428f
C169 vdd.t23 vss 0.17428f
C170 vdd.t57 vss 0.17428f
C171 vdd.t35 vss 0.17428f
C172 vdd.t41 vss 0.17428f
C173 vdd.t25 vss 0.17428f
C174 vdd.t33 vss 0.17428f
C175 vdd.t21 vss 0.17428f
C176 vdd.t49 vss 0.13071f
C177 vdd.n47 vss 0.114488f
C178 vdd.n48 vss 0.114488f
C179 vdd.n49 vss 0.08714f
C180 vdd.n50 vss 0.114488f
C181 vdd.n51 vss 0.07041f
C182 vdd.n52 vss 0.068634f
C183 vdd.n53 vss 0.2704f
C184 vdd.n54 vss 0.21187f
C185 vdd.t26 vss 0.005014f
C186 vdd.t42 vss 0.005014f
C187 vdd.n55 vss 0.010787f
C188 vdd.t16 vss 0.005014f
C189 vdd.t65 vss 0.005014f
C190 vdd.n56 vss 0.010772f
C191 vdd.t36 vss 0.005014f
C192 vdd.t58 vss 0.005014f
C193 vdd.n57 vss 0.01078f
C194 vdd.t24 vss 0.005014f
C195 vdd.t20 vss 0.005014f
C196 vdd.n58 vss 0.010776f
C197 vdd.n59 vss 0.150396f
C198 vdd.t32 vss 0.018904f
C199 vdd.n60 vss 0.181286f
C200 vdd.n61 vss 0.35924f
C201 vdd.n62 vss 0.049792f
C202 vdd.n63 vss 0.164475f
C203 vdd.n64 vss 0.028491f
C204 vdd.n65 vss 0.113062f
C205 vdd.n66 vss 0.142172f
C206 vdd.n67 vss 0.125259f
C207 vdd.n68 vss 0.12327f
C208 vdd.n69 vss 0.206776f
C209 vdd.n70 vss 0.170828f
C210 vdd.n71 vss 0.170184f
C211 vdd.n72 vss 0.142725f
C212 vdd.n73 vss 0.168715f
C213 vdd.n74 vss 0.156133f
C214 vdd.n75 vss 0.047026f
C215 vdd.n76 vss 2.27976f
C216 vdd.n77 vss 2.04931f
C217 vdd.n78 vss 0.643664f
C218 vdd.t0 vss 0.021547f
C219 vdd.n79 vss 1.8034f
C220 out.t0 vss 17.0627f
C221 out.t1 vss 0.030747f
C222 out.n0 vss 1.69316f
C223 out.n1 vss 0.319444f
C224 out.n2 vss 8.47466f
C225 out.n3 vss 0.228588f
C226 out.t21 vss 0.004354f
C227 out.t18 vss 0.004354f
C228 out.n4 vss 0.009991f
C229 out.t15 vss 0.004354f
C230 out.t13 vss 0.004354f
C231 out.n5 vss 0.009944f
C232 out.n6 vss 0.294111f
C233 out.t23 vss 0.015296f
C234 out.n7 vss 0.029896f
C235 out.t3 vss 0.004354f
C236 out.t19 vss 0.004354f
C237 out.n8 vss 0.009369f
C238 out.t10 vss 0.004354f
C239 out.t6 vss 0.004354f
C240 out.n9 vss 0.009307f
C241 out.t4 vss 0.004354f
C242 out.t9 vss 0.004354f
C243 out.n10 vss 0.009296f
C244 out.t25 vss 0.004354f
C245 out.t27 vss 0.004354f
C246 out.n11 vss 0.010391f
C247 out.t8 vss 0.004354f
C248 out.t7 vss 0.004354f
C249 out.n12 vss 0.009296f
C250 out.t20 vss 0.004354f
C251 out.t16 vss 0.004354f
C252 out.n13 vss 0.009296f
C253 out.t11 vss 0.004354f
C254 out.t12 vss 0.004354f
C255 out.n14 vss 0.009296f
C256 out.t22 vss 0.004354f
C257 out.t24 vss 0.004354f
C258 out.n15 vss 0.010471f
C259 out.t17 vss 0.004354f
C260 out.t2 vss 0.004354f
C261 out.n16 vss 0.009288f
C262 out.t14 vss 0.004354f
C263 out.t5 vss 0.004354f
C264 out.n17 vss 0.009288f
C265 out.t26 vss 0.004354f
C266 out.t28 vss 0.004354f
C267 out.n18 vss 0.011309f
C268 out.n19 vss 0.411658f
C269 out.n20 vss 0.143381f
C270 out.n21 vss 0.157433f
C271 out.n22 vss 0.179935f
C272 out.n23 vss 0.189695f
C273 out.n24 vss 0.915709f
C274 out.n25 vss 0.155485f
C275 out.n26 vss 0.184815f
C276 out.n27 vss 0.173542f
C277 out.n28 vss 0.143412f
C278 out.n29 vss 0.722411f
C279 out.n30 vss 0.351424f
C280 out.n31 vss 3.85203f
C281 p3_opamp_0.V1.n0 vss 1.40523f
C282 p3_opamp_0.V1.n1 vss 0.883305f
C283 p3_opamp_0.V1.t8 vss 0.215836f
C284 p3_opamp_0.V1.t16 vss 0.215719f
C285 p3_opamp_0.V1.t10 vss 0.215719f
C286 p3_opamp_0.V1.t12 vss 0.215719f
C287 p3_opamp_0.V1.t13 vss 0.215719f
C288 p3_opamp_0.V1.t9 vss 0.215719f
C289 p3_opamp_0.V1.t22 vss 0.215719f
C290 p3_opamp_0.V1.t14 vss 0.215719f
C291 p3_opamp_0.V1.t17 vss 0.215719f
C292 p3_opamp_0.V1.t21 vss 0.215719f
C293 p3_opamp_0.V1.t11 vss 0.215719f
C294 p3_opamp_0.V1.t25 vss 0.215719f
C295 p3_opamp_0.V1.t19 vss 0.215719f
C296 p3_opamp_0.V1.t23 vss 0.215719f
C297 p3_opamp_0.V1.t15 vss 0.215719f
C298 p3_opamp_0.V1.t18 vss 0.215719f
C299 p3_opamp_0.V1.t7 vss 0.215719f
C300 p3_opamp_0.V1.t20 vss 0.215838f
C301 p3_opamp_0.V1.t26 vss 0.215719f
C302 p3_opamp_0.V1.t24 vss 0.215719f
C303 p3_opamp_0.V1.t2 vss 0.017916f
C304 p3_opamp_0.V1.t3 vss 0.017916f
C305 p3_opamp_0.V1.n2 vss 0.038835f
C306 p3_opamp_0.V1.t0 vss 0.017916f
C307 p3_opamp_0.V1.t4 vss 0.017916f
C308 p3_opamp_0.V1.n3 vss 0.038818f
C309 p3_opamp_0.V1.t5 vss 0.069923f
C310 p3_opamp_0.V1.t1 vss 0.179078f
C311 p3_opamp_0.V1.t6 vss 0.066605f
C312 p3_opamp_0.V1.n4 vss 1.2521f
C313 twin_tee_0.c3_c4.t0 vss 14.727901f
C314 twin_tee_0.c3_c4.t2 vss 20.902302f
C315 twin_tee_0.c3_c4.n0 vss 6.25399f
C316 twin_tee_0.c3_c4.t1 vss 0.079662f
C317 p3_opamp_0.VBIAS.t0 vss 0.033592f
C318 p3_opamp_0.VBIAS.t2 vss 0.001609f
C319 p3_opamp_0.VBIAS.t8 vss 0.001609f
C320 p3_opamp_0.VBIAS.n0 vss 0.00353f
C321 p3_opamp_0.VBIAS.t6 vss 0.001609f
C322 p3_opamp_0.VBIAS.t4 vss 0.001609f
C323 p3_opamp_0.VBIAS.n1 vss 0.00353f
C324 p3_opamp_0.VBIAS.t18 vss 0.067433f
C325 p3_opamp_0.VBIAS.t16 vss 0.066149f
C326 p3_opamp_0.VBIAS.n2 vss 0.148179f
C327 p3_opamp_0.VBIAS.t14 vss 0.066149f
C328 p3_opamp_0.VBIAS.n3 vss 0.077179f
C329 p3_opamp_0.VBIAS.t19 vss 0.066149f
C330 p3_opamp_0.VBIAS.n4 vss 0.076984f
C331 p3_opamp_0.VBIAS.t17 vss 0.066149f
C332 p3_opamp_0.VBIAS.n5 vss 0.077373f
C333 p3_opamp_0.VBIAS.t15 vss 0.066149f
C334 p3_opamp_0.VBIAS.n6 vss 0.073605f
C335 p3_opamp_0.VBIAS.t13 vss 0.066286f
C336 p3_opamp_0.VBIAS.n7 vss 0.412165f
C337 p3_opamp_0.VBIAS.t12 vss 0.067681f
C338 p3_opamp_0.VBIAS.t9 vss 0.066142f
C339 p3_opamp_0.VBIAS.n8 vss 0.142758f
C340 p3_opamp_0.VBIAS.t10 vss 0.066142f
C341 p3_opamp_0.VBIAS.n9 vss 0.07339f
C342 p3_opamp_0.VBIAS.t11 vss 0.066142f
C343 p3_opamp_0.VBIAS.n10 vss 0.078801f
C344 p3_opamp_0.VBIAS.t3 vss 0.066241f
C345 p3_opamp_0.VBIAS.n11 vss 0.119554f
C346 p3_opamp_0.VBIAS.n12 vss 0.160208f
C347 p3_opamp_0.VBIAS.n13 vss 0.017329f
C348 p3_opamp_0.VBIAS.t5 vss 0.066241f
C349 p3_opamp_0.VBIAS.n14 vss 0.109887f
C350 p3_opamp_0.VBIAS.t7 vss 0.066241f
C351 p3_opamp_0.VBIAS.n15 vss 0.109887f
C352 p3_opamp_0.VBIAS.n16 vss 0.022864f
C353 p3_opamp_0.VBIAS.t1 vss 0.066241f
C354 p3_opamp_0.VBIAS.n17 vss 0.113577f
.ends

