magic
tech sky130A
magscale 1 2
timestamp 1715688618
<< psubdiff >>
rect -456 3854 2 3878
rect -456 3292 2 3316
<< psubdiffcont >>
rect -456 3316 2 3854
<< locali >>
rect -456 3854 2 3870
rect -456 3300 2 3316
<< viali >>
rect 968 4988 1438 5090
rect 4704 5004 5176 5108
rect 2538 4320 3010 4422
rect 6268 4342 6746 4446
rect -456 3376 2 3774
rect 1410 -3678 1858 -3584
rect 6446 -3678 6892 -3590
<< metal1 >>
rect -768 5116 -314 5298
rect 7806 5163 8260 5434
rect -768 5090 1460 5116
rect -768 4988 968 5090
rect 1438 4988 1460 5090
rect -768 4968 1460 4988
rect 3450 5108 5236 5122
rect 3450 5004 4704 5108
rect 5176 5004 5236 5108
rect 3450 4986 5236 5004
rect 7323 5037 8260 5163
rect -768 4796 -314 4968
rect 376 3938 524 4968
rect 3450 4436 3586 4986
rect 7323 4458 7449 5037
rect 7778 4932 8260 5037
rect 6254 4446 7454 4458
rect 2504 4422 3766 4436
rect 2504 4320 2538 4422
rect 3010 4320 3766 4422
rect 2504 4300 3766 4320
rect 3902 4300 3908 4436
rect 6254 4342 6268 4446
rect 6746 4342 7454 4446
rect 6254 4332 7454 4342
rect 7778 3952 7967 4932
rect -486 3774 42 3854
rect 376 3790 1988 3938
rect -486 3376 -456 3774
rect 2 3376 42 3774
rect -486 3242 42 3376
rect -660 2760 42 3242
rect -660 2740 -206 2760
rect -562 409 -324 2740
rect -562 171 697 409
rect 935 171 941 409
rect -562 -3556 -324 171
rect -216 170 400 171
rect 1842 106 1986 3790
rect 7762 3184 7982 3952
rect 7756 2964 7762 3184
rect 7982 2964 7988 3184
rect 836 -38 842 106
rect 986 -38 1986 106
rect 3822 -2120 3978 -2114
rect 3822 -3184 3978 -2276
rect 3822 -3340 7530 -3184
rect -562 -3584 1883 -3556
rect 7374 -3564 7530 -3340
rect -562 -3678 1410 -3584
rect 1858 -3678 1883 -3584
rect -562 -3707 1883 -3678
rect 6420 -3590 7530 -3564
rect 6420 -3678 6446 -3590
rect 6892 -3678 7530 -3590
rect -562 -3751 -324 -3707
rect 6420 -3720 7530 -3678
<< via1 >>
rect 3766 4300 3902 4436
rect 697 171 935 409
rect 7762 2964 7982 3184
rect 842 -38 986 106
rect 3822 -2276 3978 -2120
<< metal2 >>
rect 3766 4436 3902 4442
rect 3766 4220 3902 4300
rect 3766 4075 3902 4084
rect 7762 3184 7982 3190
rect 7762 2481 7982 2964
rect 7758 2271 7767 2481
rect 7977 2271 7986 2481
rect 7762 2266 7982 2271
rect 697 409 935 415
rect 935 171 1065 409
rect 1303 171 1312 409
rect 697 165 935 171
rect 842 106 986 112
rect 77 -38 86 106
rect 230 -38 842 106
rect 842 -44 986 -38
rect 3822 -1720 3978 -1711
rect 3822 -2120 3978 -1876
rect 3816 -2276 3822 -2120
rect 3978 -2276 3984 -2120
<< via2 >>
rect 3766 4084 3902 4220
rect 7767 2271 7977 2481
rect 1065 171 1303 409
rect 86 -38 230 106
rect 3822 -1876 3978 -1720
<< metal3 >>
rect 3761 4220 3907 4225
rect 3761 4084 3766 4220
rect 3902 4084 3907 4220
rect 3761 4079 3907 4084
rect 3766 4062 3902 4079
rect 3766 3920 3902 3926
rect 7762 2481 7982 2486
rect 7762 2271 7767 2481
rect 7977 2271 7982 2481
rect 1060 409 1308 414
rect 1060 171 1065 409
rect 1303 171 1373 409
rect 1611 171 1617 409
rect 1060 166 1308 171
rect 7762 159 7982 2271
rect 81 106 235 111
rect 81 -38 86 106
rect 230 -38 235 106
rect 81 -43 235 -38
rect 86 -320 230 -43
rect 7757 -59 7763 159
rect 7981 -59 7987 159
rect 7762 -60 7982 -59
rect 86 -470 230 -464
rect 3822 -1402 3978 -1396
rect 3822 -1715 3978 -1558
rect 3817 -1720 3983 -1715
rect 3817 -1876 3822 -1720
rect 3978 -1876 3983 -1720
rect 3817 -1881 3983 -1876
<< via3 >>
rect 3766 3926 3902 4062
rect 1373 171 1611 409
rect 7763 -59 7981 159
rect 86 -464 230 -320
rect 3822 -1558 3978 -1402
<< metal4 >>
rect 3765 4062 3903 4063
rect 3765 3964 3766 4062
rect 3542 3926 3766 3964
rect 3902 3964 3903 4062
rect 3902 3926 7536 3964
rect 3542 3728 7536 3926
rect 3542 2560 3778 3728
rect 7300 2448 7536 3728
rect 1716 417 1942 1932
rect 5715 417 5941 2223
rect 1372 409 1612 410
rect 1716 409 5941 417
rect 1372 171 1373 409
rect 1611 191 5941 409
rect 1611 171 1901 191
rect 1372 170 1612 171
rect 7334 159 7982 160
rect 7334 -59 7763 159
rect 7981 -59 7982 159
rect 7334 -60 7982 -59
rect 85 -320 231 -319
rect 85 -464 86 -320
rect 230 -464 231 -320
rect 85 -465 231 -464
rect 86 -570 230 -465
rect 86 -714 814 -570
rect 3564 -1158 4616 -196
rect 7334 -1028 7554 -60
rect 3822 -1401 3978 -1158
rect 3821 -1402 3979 -1401
rect 3821 -1558 3822 -1402
rect 3978 -1558 3979 -1402
rect 3821 -1559 3979 -1558
use sky130_fd_pr__res_high_po_0p35_EMSEB3  sky130_fd_pr__res_high_po_0p35_EMSEB3_0
timestamp 1715688561
transform 0 1 1978 -1 0 4711
box -533 -1246 533 1246
use sky130_fd_pr__res_high_po_0p35_EMSEB3  sky130_fd_pr__res_high_po_0p35_EMSEB3_2
timestamp 1715688561
transform 0 1 5736 -1 0 4723
box -533 -1246 533 1246
use sky130_fd_pr__cap_mim_m3_1_MRZGNS  XC1
timestamp 1715687893
transform 1 0 2035 0 1 2087
box -1686 -1540 1686 1540
use sky130_fd_pr__cap_mim_m3_1_MRZGNS  XC2
timestamp 1715687893
transform 1 0 5784 0 1 2050
box -1686 -1540 1686 1540
use sky130_fd_pr__cap_mim_m3_1_MRZGNS  XC3
timestamp 1715687893
transform 1 0 2026 0 1 -1632
box -1686 -1540 1686 1540
use sky130_fd_pr__cap_mim_m3_1_MRZGNS  XC4
timestamp 1715687893
transform 1 0 5818 0 1 -1592
box -1686 -1540 1686 1540
use sky130_fd_pr__res_high_po_0p35_4P6F7P  XR6
timestamp 1715687893
transform 0 1 4154 -1 0 -3637
box -201 -2898 201 2898
<< labels >>
flabel metal1 -616 2860 -416 3060 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 -626 5012 -426 5212 0 FreeSans 256 0 0 0 in
port 3 nsew
flabel metal1 3450 4986 4704 5122 0 FreeSans 1600 0 0 0 c1_c2
flabel metal1 7902 5004 8102 5204 0 FreeSans 256 0 0 0 out
port 2 nsew
flabel metal4 3564 -1158 4616 -196 0 FreeSans 1600 0 0 0 c3_c4
<< end >>
