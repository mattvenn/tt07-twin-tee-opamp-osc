magic
tech sky130A
magscale 1 2
timestamp 1715774553
<< viali >>
rect 4077 11305 4111 11339
rect 6101 11305 6135 11339
rect 6469 11305 6503 11339
rect 2697 11237 2731 11271
rect 6745 11237 6779 11271
rect 6961 11237 6995 11271
rect 2329 11169 2363 11203
rect 3525 11169 3559 11203
rect 3893 11169 3927 11203
rect 4261 11169 4295 11203
rect 5181 11169 5215 11203
rect 6285 11169 6319 11203
rect 6653 11169 6687 11203
rect 7481 11169 7515 11203
rect 7573 11169 7607 11203
rect 7757 11169 7791 11203
rect 8033 11169 8067 11203
rect 8401 11169 8435 11203
rect 8668 11169 8702 11203
rect 3433 11101 3467 11135
rect 3617 11101 3651 11135
rect 3709 11101 3743 11135
rect 4905 11101 4939 11135
rect 5457 11101 5491 11135
rect 7205 11101 7239 11135
rect 7389 11101 7423 11135
rect 8217 11101 8251 11135
rect 10425 11101 10459 11135
rect 10793 11101 10827 11135
rect 3249 11033 3283 11067
rect 5365 11033 5399 11067
rect 7113 11033 7147 11067
rect 7481 11033 7515 11067
rect 2697 10965 2731 10999
rect 2881 10965 2915 10999
rect 4997 10965 5031 10999
rect 6929 10965 6963 10999
rect 7573 10965 7607 10999
rect 7849 10965 7883 10999
rect 9781 10965 9815 10999
rect 9873 10965 9907 10999
rect 1317 10761 1351 10795
rect 1685 10761 1719 10795
rect 2881 10761 2915 10795
rect 3525 10693 3559 10727
rect 6653 10693 6687 10727
rect 8217 10693 8251 10727
rect 1961 10625 1995 10659
rect 3893 10625 3927 10659
rect 4813 10625 4847 10659
rect 7849 10625 7883 10659
rect 8953 10625 8987 10659
rect 10793 10625 10827 10659
rect 1501 10557 1535 10591
rect 1869 10557 1903 10591
rect 3065 10557 3099 10591
rect 3249 10557 3283 10591
rect 3341 10557 3375 10591
rect 3801 10557 3835 10591
rect 3985 10557 4019 10591
rect 4077 10557 4111 10591
rect 5181 10557 5215 10591
rect 5273 10557 5307 10591
rect 7389 10557 7423 10591
rect 7665 10557 7699 10591
rect 7941 10557 7975 10591
rect 11069 10557 11103 10591
rect 3525 10489 3559 10523
rect 4261 10489 4295 10523
rect 5518 10489 5552 10523
rect 8217 10489 8251 10523
rect 8401 10489 8435 10523
rect 2605 10421 2639 10455
rect 3617 10421 3651 10455
rect 5089 10421 5123 10455
rect 6745 10421 6779 10455
rect 7481 10421 7515 10455
rect 8033 10421 8067 10455
rect 9321 10421 9355 10455
rect 3249 10217 3283 10251
rect 5181 10217 5215 10251
rect 8585 10217 8619 10251
rect 9505 10217 9539 10251
rect 1409 10149 1443 10183
rect 4568 10149 4602 10183
rect 1041 10081 1075 10115
rect 1225 10081 1259 10115
rect 1317 10081 1351 10115
rect 1593 10081 1627 10115
rect 2798 10081 2832 10115
rect 3157 10081 3191 10115
rect 3341 10081 3375 10115
rect 4905 10081 4939 10115
rect 5089 10081 5123 10115
rect 5365 10081 5399 10115
rect 5549 10081 5583 10115
rect 5641 10081 5675 10115
rect 6009 10081 6043 10115
rect 7021 10081 7055 10115
rect 7113 10081 7147 10115
rect 7380 10081 7414 10115
rect 9137 10081 9171 10115
rect 9321 10081 9355 10115
rect 10609 10081 10643 10115
rect 10793 10081 10827 10115
rect 3065 10013 3099 10047
rect 4813 10013 4847 10047
rect 4997 10013 5031 10047
rect 6285 10013 6319 10047
rect 6377 10013 6411 10047
rect 10241 10013 10275 10047
rect 10517 10013 10551 10047
rect 1685 9945 1719 9979
rect 6193 9945 6227 9979
rect 1225 9877 1259 9911
rect 1593 9877 1627 9911
rect 3433 9877 3467 9911
rect 5825 9877 5859 9911
rect 8493 9877 8527 9911
rect 10609 9877 10643 9911
rect 1317 9673 1351 9707
rect 5273 9673 5307 9707
rect 7021 9673 7055 9707
rect 7941 9673 7975 9707
rect 8861 9673 8895 9707
rect 1133 9605 1167 9639
rect 2881 9605 2915 9639
rect 4997 9605 5031 9639
rect 7665 9605 7699 9639
rect 8493 9605 8527 9639
rect 10333 9605 10367 9639
rect 2697 9537 2731 9571
rect 5641 9537 5675 9571
rect 10977 9537 11011 9571
rect 1225 9469 1259 9503
rect 2430 9469 2464 9503
rect 3065 9469 3099 9503
rect 3433 9469 3467 9503
rect 5181 9469 5215 9503
rect 5549 9469 5583 9503
rect 7389 9469 7423 9503
rect 8401 9469 8435 9503
rect 8677 9469 8711 9503
rect 8953 9469 8987 9503
rect 3678 9401 3712 9435
rect 5273 9401 5307 9435
rect 5908 9401 5942 9435
rect 7481 9401 7515 9435
rect 8125 9401 8159 9435
rect 9198 9401 9232 9435
rect 4813 9333 4847 9367
rect 5457 9333 5491 9367
rect 7113 9333 7147 9367
rect 7297 9333 7331 9367
rect 7757 9333 7791 9367
rect 7925 9333 7959 9367
rect 10425 9333 10459 9367
rect 2421 9129 2455 9163
rect 3249 9129 3283 9163
rect 3417 9129 3451 9163
rect 5825 9129 5859 9163
rect 6561 9129 6595 9163
rect 8033 9129 8067 9163
rect 3617 9061 3651 9095
rect 5457 9061 5491 9095
rect 8585 9061 8619 9095
rect 10333 9061 10367 9095
rect 2605 8993 2639 9027
rect 2881 8993 2915 9027
rect 6009 8993 6043 9027
rect 7849 8993 7883 9027
rect 8217 8993 8251 9027
rect 8493 8993 8527 9027
rect 10609 8993 10643 9027
rect 2697 8925 2731 8959
rect 2789 8925 2823 8959
rect 3709 8925 3743 8959
rect 10793 8925 10827 8959
rect 3433 8789 3467 8823
rect 8401 8789 8435 8823
rect 10425 8789 10459 8823
rect 2881 8585 2915 8619
rect 4261 8585 4295 8619
rect 7481 8585 7515 8619
rect 8769 8585 8803 8619
rect 3433 8517 3467 8551
rect 4169 8517 4203 8551
rect 6377 8517 6411 8551
rect 8125 8517 8159 8551
rect 5641 8449 5675 8483
rect 3065 8381 3099 8415
rect 3249 8381 3283 8415
rect 3433 8381 3467 8415
rect 3525 8381 3559 8415
rect 3709 8381 3743 8415
rect 3801 8381 3835 8415
rect 3893 8381 3927 8415
rect 3985 8381 4019 8415
rect 4905 8381 4939 8415
rect 5549 8381 5583 8415
rect 5825 8381 5859 8415
rect 6193 8381 6227 8415
rect 6469 8381 6503 8415
rect 6745 8381 6779 8415
rect 6837 8381 6871 8415
rect 6929 8381 6963 8415
rect 7205 8381 7239 8415
rect 7297 8381 7331 8415
rect 7941 8381 7975 8415
rect 8217 8381 8251 8415
rect 8585 8381 8619 8415
rect 8861 8381 8895 8415
rect 8953 8381 8987 8415
rect 10977 8381 11011 8415
rect 4169 8313 4203 8347
rect 4997 8313 5031 8347
rect 5365 8313 5399 8347
rect 6561 8313 6595 8347
rect 8401 8313 8435 8347
rect 9198 8313 9232 8347
rect 10425 8313 10459 8347
rect 3801 8245 3835 8279
rect 5181 8245 5215 8279
rect 5273 8245 5307 8279
rect 6009 8245 6043 8279
rect 7757 8245 7791 8279
rect 10333 8245 10367 8279
rect 4813 8041 4847 8075
rect 6745 8041 6779 8075
rect 7481 8041 7515 8075
rect 8401 8041 8435 8075
rect 8953 8041 8987 8075
rect 10241 8041 10275 8075
rect 10609 8041 10643 8075
rect 8493 7973 8527 8007
rect 10425 7973 10459 8007
rect 2789 7905 2823 7939
rect 3065 7905 3099 7939
rect 3157 7905 3191 7939
rect 3424 7905 3458 7939
rect 6377 7905 6411 7939
rect 7757 7905 7791 7939
rect 7849 7905 7883 7939
rect 8125 7905 8159 7939
rect 8309 7905 8343 7939
rect 9873 7905 9907 7939
rect 10057 7905 10091 7939
rect 10517 7905 10551 7939
rect 5457 7837 5491 7871
rect 7389 7837 7423 7871
rect 7665 7837 7699 7871
rect 7941 7837 7975 7871
rect 9505 7837 9539 7871
rect 10149 7837 10183 7871
rect 10793 7769 10827 7803
rect 2605 7701 2639 7735
rect 2973 7701 3007 7735
rect 4537 7701 4571 7735
rect 5825 7701 5859 7735
rect 8677 7701 8711 7735
rect 9689 7701 9723 7735
rect 2421 7497 2455 7531
rect 3433 7497 3467 7531
rect 5457 7497 5491 7531
rect 7021 7497 7055 7531
rect 7389 7497 7423 7531
rect 8217 7497 8251 7531
rect 9321 7497 9355 7531
rect 1777 7361 1811 7395
rect 3065 7361 3099 7395
rect 9229 7361 9263 7395
rect 10241 7361 10275 7395
rect 3709 7293 3743 7327
rect 3965 7293 3999 7327
rect 5181 7293 5215 7327
rect 5457 7293 5491 7327
rect 5641 7293 5675 7327
rect 5908 7293 5942 7327
rect 7113 7293 7147 7327
rect 7665 7293 7699 7327
rect 8953 7293 8987 7327
rect 9321 7293 9355 7327
rect 9505 7293 9539 7327
rect 10425 7293 10459 7327
rect 2329 7225 2363 7259
rect 3249 7225 3283 7259
rect 3465 7225 3499 7259
rect 7389 7225 7423 7259
rect 3617 7157 3651 7191
rect 5089 7157 5123 7191
rect 5273 7157 5307 7191
rect 7205 7157 7239 7191
rect 9597 7157 9631 7191
rect 10977 7157 11011 7191
rect 3617 6953 3651 6987
rect 9229 6953 9263 6987
rect 10701 6953 10735 6987
rect 2237 6817 2271 6851
rect 2504 6817 2538 6851
rect 3976 6817 4010 6851
rect 5181 6817 5215 6851
rect 5365 6817 5399 6851
rect 6101 6817 6135 6851
rect 6285 6817 6319 6851
rect 6644 6817 6678 6851
rect 8116 6817 8150 6851
rect 9588 6817 9622 6851
rect 3709 6749 3743 6783
rect 6377 6749 6411 6783
rect 7849 6749 7883 6783
rect 9321 6749 9355 6783
rect 5089 6681 5123 6715
rect 6285 6681 6319 6715
rect 5365 6613 5399 6647
rect 7757 6613 7791 6647
rect 3709 6409 3743 6443
rect 4169 6409 4203 6443
rect 8125 6409 8159 6443
rect 8953 6409 8987 6443
rect 9505 6409 9539 6443
rect 4537 6341 4571 6375
rect 7205 6341 7239 6375
rect 8677 6341 8711 6375
rect 5825 6273 5859 6307
rect 7573 6273 7607 6307
rect 9413 6273 9447 6307
rect 3985 6205 4019 6239
rect 4353 6205 4387 6239
rect 4629 6205 4663 6239
rect 4905 6205 4939 6239
rect 5457 6205 5491 6239
rect 6092 6205 6126 6239
rect 8861 6205 8895 6239
rect 9137 6205 9171 6239
rect 9321 6205 9355 6239
rect 10885 6205 10919 6239
rect 3709 6137 3743 6171
rect 10640 6137 10674 6171
rect 3893 6069 3927 6103
rect 7665 5865 7699 5899
rect 8769 5865 8803 5899
rect 9229 5865 9263 5899
rect 10701 5865 10735 5899
rect 7389 5729 7423 5763
rect 7481 5729 7515 5763
rect 8677 5729 8711 5763
rect 8861 5729 8895 5763
rect 9137 5729 9171 5763
rect 9413 5729 9447 5763
rect 9873 5729 9907 5763
rect 10425 5729 10459 5763
rect 10517 5729 10551 5763
rect 10793 5729 10827 5763
rect 9413 5593 9447 5627
rect 10517 5593 10551 5627
rect 10333 5321 10367 5355
rect 10609 5321 10643 5355
rect 10425 5253 10459 5287
rect 9965 5185 9999 5219
rect 10149 5117 10183 5151
rect 10577 5049 10611 5083
rect 10793 5049 10827 5083
rect 10793 4777 10827 4811
rect 10517 4641 10551 4675
rect 10701 4641 10735 4675
rect 10793 4641 10827 4675
<< metal1 >>
rect 3970 11636 3976 11688
rect 4028 11676 4034 11688
rect 7834 11676 7840 11688
rect 4028 11648 7840 11676
rect 4028 11636 4034 11648
rect 7834 11636 7840 11648
rect 7892 11676 7898 11688
rect 9582 11676 9588 11688
rect 7892 11648 9588 11676
rect 7892 11636 7898 11648
rect 9582 11636 9588 11648
rect 9640 11636 9646 11688
rect 6638 11568 6644 11620
rect 6696 11608 6702 11620
rect 8018 11608 8024 11620
rect 6696 11580 8024 11608
rect 6696 11568 6702 11580
rect 8018 11568 8024 11580
rect 8076 11568 8082 11620
rect 8294 11568 8300 11620
rect 8352 11608 8358 11620
rect 8478 11608 8484 11620
rect 8352 11580 8484 11608
rect 8352 11568 8358 11580
rect 8478 11568 8484 11580
rect 8536 11568 8542 11620
rect 2866 11500 2872 11552
rect 2924 11540 2930 11552
rect 3326 11540 3332 11552
rect 2924 11512 3332 11540
rect 2924 11500 2930 11512
rect 3326 11500 3332 11512
rect 3384 11500 3390 11552
rect 5902 11500 5908 11552
rect 5960 11540 5966 11552
rect 6178 11540 6184 11552
rect 5960 11512 6184 11540
rect 5960 11500 5966 11512
rect 6178 11500 6184 11512
rect 6236 11500 6242 11552
rect 7190 11500 7196 11552
rect 7248 11540 7254 11552
rect 9490 11540 9496 11552
rect 7248 11512 9496 11540
rect 7248 11500 7254 11512
rect 9490 11500 9496 11512
rect 9548 11500 9554 11552
rect 552 11450 11568 11472
rect 552 11398 3112 11450
rect 3164 11398 3176 11450
rect 3228 11398 3240 11450
rect 3292 11398 3304 11450
rect 3356 11398 3368 11450
rect 3420 11398 5826 11450
rect 5878 11398 5890 11450
rect 5942 11398 5954 11450
rect 6006 11398 6018 11450
rect 6070 11398 6082 11450
rect 6134 11398 8540 11450
rect 8592 11398 8604 11450
rect 8656 11398 8668 11450
rect 8720 11398 8732 11450
rect 8784 11398 8796 11450
rect 8848 11398 11254 11450
rect 11306 11398 11318 11450
rect 11370 11398 11382 11450
rect 11434 11398 11446 11450
rect 11498 11398 11510 11450
rect 11562 11398 11568 11450
rect 552 11376 11568 11398
rect 4065 11339 4123 11345
rect 4065 11305 4077 11339
rect 4111 11336 4123 11339
rect 4614 11336 4620 11348
rect 4111 11308 4620 11336
rect 4111 11305 4123 11308
rect 4065 11299 4123 11305
rect 4614 11296 4620 11308
rect 4672 11296 4678 11348
rect 6089 11339 6147 11345
rect 6089 11305 6101 11339
rect 6135 11336 6147 11339
rect 6178 11336 6184 11348
rect 6135 11308 6184 11336
rect 6135 11305 6147 11308
rect 6089 11299 6147 11305
rect 6178 11296 6184 11308
rect 6236 11296 6242 11348
rect 6457 11339 6515 11345
rect 6457 11305 6469 11339
rect 6503 11336 6515 11339
rect 8294 11336 8300 11348
rect 6503 11308 8300 11336
rect 6503 11305 6515 11308
rect 6457 11299 6515 11305
rect 8294 11296 8300 11308
rect 8352 11296 8358 11348
rect 2682 11228 2688 11280
rect 2740 11228 2746 11280
rect 3970 11268 3976 11280
rect 2976 11240 3976 11268
rect 2317 11203 2375 11209
rect 2317 11169 2329 11203
rect 2363 11200 2375 11203
rect 2976 11200 3004 11240
rect 3970 11228 3976 11240
rect 4028 11228 4034 11280
rect 6733 11271 6791 11277
rect 6733 11237 6745 11271
rect 6779 11237 6791 11271
rect 6733 11231 6791 11237
rect 6949 11271 7007 11277
rect 6949 11237 6961 11271
rect 6995 11268 7007 11271
rect 7650 11268 7656 11280
rect 6995 11240 7656 11268
rect 6995 11237 7007 11240
rect 6949 11231 7007 11237
rect 2363 11172 3004 11200
rect 2363 11169 2375 11172
rect 2317 11163 2375 11169
rect 3050 11160 3056 11212
rect 3108 11200 3114 11212
rect 3513 11203 3571 11209
rect 3513 11200 3525 11203
rect 3108 11172 3525 11200
rect 3108 11160 3114 11172
rect 3513 11169 3525 11172
rect 3559 11169 3571 11203
rect 3881 11203 3939 11209
rect 3881 11200 3893 11203
rect 3513 11163 3571 11169
rect 3620 11172 3893 11200
rect 3620 11144 3648 11172
rect 3881 11169 3893 11172
rect 3927 11200 3939 11203
rect 4249 11203 4307 11209
rect 4249 11200 4261 11203
rect 3927 11172 4261 11200
rect 3927 11169 3939 11172
rect 3881 11163 3939 11169
rect 4249 11169 4261 11172
rect 4295 11169 4307 11203
rect 4249 11163 4307 11169
rect 5166 11160 5172 11212
rect 5224 11160 5230 11212
rect 6273 11203 6331 11209
rect 6273 11169 6285 11203
rect 6319 11169 6331 11203
rect 6273 11163 6331 11169
rect 3421 11135 3479 11141
rect 3421 11101 3433 11135
rect 3467 11101 3479 11135
rect 3421 11095 3479 11101
rect 3237 11067 3295 11073
rect 3237 11064 3249 11067
rect 2700 11036 3249 11064
rect 2700 11005 2728 11036
rect 3237 11033 3249 11036
rect 3283 11033 3295 11067
rect 3436 11064 3464 11095
rect 3602 11092 3608 11144
rect 3660 11092 3666 11144
rect 3697 11135 3755 11141
rect 3697 11101 3709 11135
rect 3743 11132 3755 11135
rect 3786 11132 3792 11144
rect 3743 11104 3792 11132
rect 3743 11101 3755 11104
rect 3697 11095 3755 11101
rect 3786 11092 3792 11104
rect 3844 11092 3850 11144
rect 4893 11135 4951 11141
rect 4893 11101 4905 11135
rect 4939 11132 4951 11135
rect 5445 11135 5503 11141
rect 5445 11132 5457 11135
rect 4939 11104 5457 11132
rect 4939 11101 4951 11104
rect 4893 11095 4951 11101
rect 5445 11101 5457 11104
rect 5491 11101 5503 11135
rect 6288 11132 6316 11163
rect 6638 11160 6644 11212
rect 6696 11160 6702 11212
rect 6748 11200 6776 11231
rect 7650 11228 7656 11240
rect 7708 11228 7714 11280
rect 11054 11268 11060 11280
rect 8404 11240 11060 11268
rect 6748 11172 7052 11200
rect 7024 11144 7052 11172
rect 7098 11160 7104 11212
rect 7156 11200 7162 11212
rect 7469 11203 7527 11209
rect 7469 11200 7481 11203
rect 7156 11172 7481 11200
rect 7156 11160 7162 11172
rect 7469 11169 7481 11172
rect 7515 11169 7527 11203
rect 7469 11163 7527 11169
rect 7558 11160 7564 11212
rect 7616 11160 7622 11212
rect 7745 11203 7803 11209
rect 7745 11169 7757 11203
rect 7791 11200 7803 11203
rect 7834 11200 7840 11212
rect 7791 11172 7840 11200
rect 7791 11169 7803 11172
rect 7745 11163 7803 11169
rect 7834 11160 7840 11172
rect 7892 11160 7898 11212
rect 8018 11160 8024 11212
rect 8076 11160 8082 11212
rect 8404 11209 8432 11240
rect 11054 11228 11060 11240
rect 11112 11228 11118 11280
rect 8389 11203 8447 11209
rect 8389 11169 8401 11203
rect 8435 11169 8447 11203
rect 8389 11163 8447 11169
rect 8656 11203 8714 11209
rect 8656 11169 8668 11203
rect 8702 11200 8714 11203
rect 8938 11200 8944 11212
rect 8702 11172 8944 11200
rect 8702 11169 8714 11172
rect 8656 11163 8714 11169
rect 8938 11160 8944 11172
rect 8996 11160 9002 11212
rect 6914 11132 6920 11144
rect 6288 11104 6920 11132
rect 5445 11095 5503 11101
rect 6914 11092 6920 11104
rect 6972 11092 6978 11144
rect 7006 11092 7012 11144
rect 7064 11092 7070 11144
rect 7190 11092 7196 11144
rect 7248 11092 7254 11144
rect 7377 11135 7435 11141
rect 7377 11101 7389 11135
rect 7423 11132 7435 11135
rect 8110 11132 8116 11144
rect 7423 11104 8116 11132
rect 7423 11101 7435 11104
rect 7377 11095 7435 11101
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 8205 11135 8263 11141
rect 8205 11101 8217 11135
rect 8251 11101 8263 11135
rect 10413 11135 10471 11141
rect 10413 11132 10425 11135
rect 8205 11095 8263 11101
rect 9784 11104 10425 11132
rect 5353 11067 5411 11073
rect 5353 11064 5365 11067
rect 3436 11036 5365 11064
rect 3237 11027 3295 11033
rect 3712 11008 3740 11036
rect 5353 11033 5365 11036
rect 5399 11033 5411 11067
rect 5353 11027 5411 11033
rect 5534 11024 5540 11076
rect 5592 11064 5598 11076
rect 7101 11067 7159 11073
rect 7101 11064 7113 11067
rect 5592 11036 7113 11064
rect 5592 11024 5598 11036
rect 7101 11033 7113 11036
rect 7147 11064 7159 11067
rect 7282 11064 7288 11076
rect 7147 11036 7288 11064
rect 7147 11033 7159 11036
rect 7101 11027 7159 11033
rect 7282 11024 7288 11036
rect 7340 11024 7346 11076
rect 7469 11067 7527 11073
rect 7469 11033 7481 11067
rect 7515 11064 7527 11067
rect 7650 11064 7656 11076
rect 7515 11036 7656 11064
rect 7515 11033 7527 11036
rect 7469 11027 7527 11033
rect 7650 11024 7656 11036
rect 7708 11024 7714 11076
rect 7926 11024 7932 11076
rect 7984 11064 7990 11076
rect 8220 11064 8248 11095
rect 7984 11036 8248 11064
rect 7984 11024 7990 11036
rect 2685 10999 2743 11005
rect 2685 10965 2697 10999
rect 2731 10965 2743 10999
rect 2685 10959 2743 10965
rect 2869 10999 2927 11005
rect 2869 10965 2881 10999
rect 2915 10996 2927 10999
rect 2958 10996 2964 11008
rect 2915 10968 2964 10996
rect 2915 10965 2927 10968
rect 2869 10959 2927 10965
rect 2958 10956 2964 10968
rect 3016 10956 3022 11008
rect 3694 10956 3700 11008
rect 3752 10956 3758 11008
rect 4982 10956 4988 11008
rect 5040 10956 5046 11008
rect 6730 10956 6736 11008
rect 6788 10996 6794 11008
rect 6917 10999 6975 11005
rect 6917 10996 6929 10999
rect 6788 10968 6929 10996
rect 6788 10956 6794 10968
rect 6917 10965 6929 10968
rect 6963 10965 6975 10999
rect 6917 10959 6975 10965
rect 7558 10956 7564 11008
rect 7616 10956 7622 11008
rect 7742 10956 7748 11008
rect 7800 10996 7806 11008
rect 7837 10999 7895 11005
rect 7837 10996 7849 10999
rect 7800 10968 7849 10996
rect 7800 10956 7806 10968
rect 7837 10965 7849 10968
rect 7883 10965 7895 10999
rect 8220 10996 8248 11036
rect 9784 11005 9812 11104
rect 10413 11101 10425 11104
rect 10459 11101 10471 11135
rect 10413 11095 10471 11101
rect 10778 11092 10784 11144
rect 10836 11092 10842 11144
rect 9769 10999 9827 11005
rect 9769 10996 9781 10999
rect 8220 10968 9781 10996
rect 7837 10959 7895 10965
rect 9769 10965 9781 10968
rect 9815 10965 9827 10999
rect 9769 10959 9827 10965
rect 9861 10999 9919 11005
rect 9861 10965 9873 10999
rect 9907 10996 9919 10999
rect 10226 10996 10232 11008
rect 9907 10968 10232 10996
rect 9907 10965 9919 10968
rect 9861 10959 9919 10965
rect 10226 10956 10232 10968
rect 10284 10956 10290 11008
rect 552 10906 11408 10928
rect 552 10854 1755 10906
rect 1807 10854 1819 10906
rect 1871 10854 1883 10906
rect 1935 10854 1947 10906
rect 1999 10854 2011 10906
rect 2063 10854 4469 10906
rect 4521 10854 4533 10906
rect 4585 10854 4597 10906
rect 4649 10854 4661 10906
rect 4713 10854 4725 10906
rect 4777 10854 7183 10906
rect 7235 10854 7247 10906
rect 7299 10854 7311 10906
rect 7363 10854 7375 10906
rect 7427 10854 7439 10906
rect 7491 10854 9897 10906
rect 9949 10854 9961 10906
rect 10013 10854 10025 10906
rect 10077 10854 10089 10906
rect 10141 10854 10153 10906
rect 10205 10854 11408 10906
rect 552 10832 11408 10854
rect 750 10752 756 10804
rect 808 10792 814 10804
rect 1305 10795 1363 10801
rect 1305 10792 1317 10795
rect 808 10764 1317 10792
rect 808 10752 814 10764
rect 1305 10761 1317 10764
rect 1351 10761 1363 10795
rect 1305 10755 1363 10761
rect 1673 10795 1731 10801
rect 1673 10761 1685 10795
rect 1719 10792 1731 10795
rect 2130 10792 2136 10804
rect 1719 10764 2136 10792
rect 1719 10761 1731 10764
rect 1673 10755 1731 10761
rect 2130 10752 2136 10764
rect 2188 10752 2194 10804
rect 2866 10752 2872 10804
rect 2924 10752 2930 10804
rect 3050 10752 3056 10804
rect 3108 10792 3114 10804
rect 3108 10764 4108 10792
rect 3108 10752 3114 10764
rect 4080 10736 4108 10764
rect 6730 10752 6736 10804
rect 6788 10792 6794 10804
rect 8294 10792 8300 10804
rect 6788 10764 8300 10792
rect 6788 10752 6794 10764
rect 1026 10684 1032 10736
rect 1084 10724 1090 10736
rect 3513 10727 3571 10733
rect 3513 10724 3525 10727
rect 1084 10696 3525 10724
rect 1084 10684 1090 10696
rect 3513 10693 3525 10696
rect 3559 10693 3571 10727
rect 3513 10687 3571 10693
rect 3786 10684 3792 10736
rect 3844 10684 3850 10736
rect 4062 10684 4068 10736
rect 4120 10684 4126 10736
rect 6641 10727 6699 10733
rect 6641 10693 6653 10727
rect 6687 10724 6699 10727
rect 6914 10724 6920 10736
rect 6687 10696 6920 10724
rect 6687 10693 6699 10696
rect 6641 10687 6699 10693
rect 6914 10684 6920 10696
rect 6972 10724 6978 10736
rect 6972 10696 7420 10724
rect 6972 10684 6978 10696
rect 1949 10659 2007 10665
rect 1949 10656 1961 10659
rect 1504 10628 1961 10656
rect 1302 10548 1308 10600
rect 1360 10588 1366 10600
rect 1504 10597 1532 10628
rect 1949 10625 1961 10628
rect 1995 10625 2007 10659
rect 3804 10656 3832 10684
rect 1949 10619 2007 10625
rect 2700 10628 3832 10656
rect 3881 10659 3939 10665
rect 1489 10591 1547 10597
rect 1489 10588 1501 10591
rect 1360 10560 1501 10588
rect 1360 10548 1366 10560
rect 1489 10557 1501 10560
rect 1535 10557 1547 10591
rect 1489 10551 1547 10557
rect 1670 10548 1676 10600
rect 1728 10588 1734 10600
rect 1857 10591 1915 10597
rect 1857 10588 1869 10591
rect 1728 10560 1869 10588
rect 1728 10548 1734 10560
rect 1857 10557 1869 10560
rect 1903 10588 1915 10591
rect 2700 10588 2728 10628
rect 3881 10625 3893 10659
rect 3927 10656 3939 10659
rect 4080 10656 4108 10684
rect 4801 10659 4859 10665
rect 4801 10656 4813 10659
rect 3927 10628 4813 10656
rect 3927 10625 3939 10628
rect 3881 10619 3939 10625
rect 4801 10625 4813 10628
rect 4847 10625 4859 10659
rect 4801 10619 4859 10625
rect 5184 10628 5396 10656
rect 1903 10560 2728 10588
rect 1903 10557 1915 10560
rect 1857 10551 1915 10557
rect 3050 10548 3056 10600
rect 3108 10548 3114 10600
rect 3234 10548 3240 10600
rect 3292 10548 3298 10600
rect 3329 10591 3387 10597
rect 3329 10557 3341 10591
rect 3375 10588 3387 10591
rect 3602 10588 3608 10600
rect 3375 10560 3608 10588
rect 3375 10557 3387 10560
rect 3329 10551 3387 10557
rect 3602 10548 3608 10560
rect 3660 10548 3666 10600
rect 3694 10548 3700 10600
rect 3752 10588 3758 10600
rect 3789 10591 3847 10597
rect 3789 10588 3801 10591
rect 3752 10560 3801 10588
rect 3752 10548 3758 10560
rect 3789 10557 3801 10560
rect 3835 10557 3847 10591
rect 3789 10551 3847 10557
rect 3970 10548 3976 10600
rect 4028 10548 4034 10600
rect 4065 10591 4123 10597
rect 4065 10557 4077 10591
rect 4111 10588 4123 10591
rect 4154 10588 4160 10600
rect 4111 10560 4160 10588
rect 4111 10557 4123 10560
rect 4065 10551 4123 10557
rect 4154 10548 4160 10560
rect 4212 10548 4218 10600
rect 5184 10597 5212 10628
rect 5169 10591 5227 10597
rect 5169 10557 5181 10591
rect 5215 10557 5227 10591
rect 5169 10551 5227 10557
rect 5261 10591 5319 10597
rect 5261 10557 5273 10591
rect 5307 10557 5319 10591
rect 5368 10588 5396 10628
rect 7392 10597 7420 10696
rect 7852 10665 7880 10764
rect 8294 10752 8300 10764
rect 8352 10752 8358 10804
rect 8202 10684 8208 10736
rect 8260 10684 8266 10736
rect 7837 10659 7895 10665
rect 7837 10625 7849 10659
rect 7883 10625 7895 10659
rect 7837 10619 7895 10625
rect 7377 10591 7435 10597
rect 5368 10560 5764 10588
rect 5261 10551 5319 10557
rect 1210 10480 1216 10532
rect 1268 10520 1274 10532
rect 3513 10523 3571 10529
rect 1268 10492 3464 10520
rect 1268 10480 1274 10492
rect 2590 10412 2596 10464
rect 2648 10412 2654 10464
rect 3436 10452 3464 10492
rect 3513 10489 3525 10523
rect 3559 10520 3571 10523
rect 4249 10523 4307 10529
rect 4249 10520 4261 10523
rect 3559 10492 4261 10520
rect 3559 10489 3571 10492
rect 3513 10483 3571 10489
rect 4249 10489 4261 10492
rect 4295 10489 4307 10523
rect 4249 10483 4307 10489
rect 4798 10480 4804 10532
rect 4856 10520 4862 10532
rect 5276 10520 5304 10551
rect 5736 10532 5764 10560
rect 7377 10557 7389 10591
rect 7423 10588 7435 10591
rect 7466 10588 7472 10600
rect 7423 10560 7472 10588
rect 7423 10557 7435 10560
rect 7377 10551 7435 10557
rect 7466 10548 7472 10560
rect 7524 10548 7530 10600
rect 7653 10591 7711 10597
rect 7653 10557 7665 10591
rect 7699 10588 7711 10591
rect 7742 10588 7748 10600
rect 7699 10560 7748 10588
rect 7699 10557 7711 10560
rect 7653 10551 7711 10557
rect 7742 10548 7748 10560
rect 7800 10548 7806 10600
rect 7852 10588 7880 10619
rect 8018 10616 8024 10668
rect 8076 10656 8082 10668
rect 8941 10659 8999 10665
rect 8941 10656 8953 10659
rect 8076 10628 8953 10656
rect 8076 10616 8082 10628
rect 8941 10625 8953 10628
rect 8987 10625 8999 10659
rect 8941 10619 8999 10625
rect 10778 10616 10784 10668
rect 10836 10616 10842 10668
rect 7929 10591 7987 10597
rect 7929 10588 7941 10591
rect 7852 10560 7941 10588
rect 7929 10557 7941 10560
rect 7975 10557 7987 10591
rect 7929 10551 7987 10557
rect 8036 10560 8524 10588
rect 4856 10492 5304 10520
rect 4856 10480 4862 10492
rect 5350 10480 5356 10532
rect 5408 10520 5414 10532
rect 5506 10523 5564 10529
rect 5506 10520 5518 10523
rect 5408 10492 5518 10520
rect 5408 10480 5414 10492
rect 5506 10489 5518 10492
rect 5552 10489 5564 10523
rect 5506 10483 5564 10489
rect 5718 10480 5724 10532
rect 5776 10480 5782 10532
rect 8036 10520 8064 10560
rect 6564 10492 8064 10520
rect 8205 10523 8263 10529
rect 3605 10455 3663 10461
rect 3605 10452 3617 10455
rect 3436 10424 3617 10452
rect 3605 10421 3617 10424
rect 3651 10421 3663 10455
rect 3605 10415 3663 10421
rect 5077 10455 5135 10461
rect 5077 10421 5089 10455
rect 5123 10452 5135 10455
rect 6564 10452 6592 10492
rect 8205 10489 8217 10523
rect 8251 10520 8263 10523
rect 8389 10523 8447 10529
rect 8389 10520 8401 10523
rect 8251 10492 8401 10520
rect 8251 10489 8263 10492
rect 8205 10483 8263 10489
rect 8389 10489 8401 10492
rect 8435 10489 8447 10523
rect 8496 10520 8524 10560
rect 11054 10548 11060 10600
rect 11112 10548 11118 10600
rect 8496 10492 9614 10520
rect 8389 10483 8447 10489
rect 5123 10424 6592 10452
rect 5123 10421 5135 10424
rect 5077 10415 5135 10421
rect 6730 10412 6736 10464
rect 6788 10412 6794 10464
rect 7098 10412 7104 10464
rect 7156 10452 7162 10464
rect 7469 10455 7527 10461
rect 7469 10452 7481 10455
rect 7156 10424 7481 10452
rect 7156 10412 7162 10424
rect 7469 10421 7481 10424
rect 7515 10421 7527 10455
rect 7469 10415 7527 10421
rect 7926 10412 7932 10464
rect 7984 10452 7990 10464
rect 8021 10455 8079 10461
rect 8021 10452 8033 10455
rect 7984 10424 8033 10452
rect 7984 10412 7990 10424
rect 8021 10421 8033 10424
rect 8067 10421 8079 10455
rect 8021 10415 8079 10421
rect 9306 10412 9312 10464
rect 9364 10412 9370 10464
rect 552 10362 11568 10384
rect 552 10310 3112 10362
rect 3164 10310 3176 10362
rect 3228 10310 3240 10362
rect 3292 10310 3304 10362
rect 3356 10310 3368 10362
rect 3420 10310 5826 10362
rect 5878 10310 5890 10362
rect 5942 10310 5954 10362
rect 6006 10310 6018 10362
rect 6070 10310 6082 10362
rect 6134 10310 8540 10362
rect 8592 10310 8604 10362
rect 8656 10310 8668 10362
rect 8720 10310 8732 10362
rect 8784 10310 8796 10362
rect 8848 10310 11254 10362
rect 11306 10310 11318 10362
rect 11370 10310 11382 10362
rect 11434 10310 11446 10362
rect 11498 10310 11510 10362
rect 11562 10310 11568 10362
rect 552 10288 11568 10310
rect 2682 10248 2688 10260
rect 1504 10220 2688 10248
rect 1118 10140 1124 10192
rect 1176 10180 1182 10192
rect 1397 10183 1455 10189
rect 1397 10180 1409 10183
rect 1176 10152 1409 10180
rect 1176 10140 1182 10152
rect 1397 10149 1409 10152
rect 1443 10149 1455 10183
rect 1397 10143 1455 10149
rect 1026 10072 1032 10124
rect 1084 10072 1090 10124
rect 1210 10072 1216 10124
rect 1268 10072 1274 10124
rect 1305 10115 1363 10121
rect 1305 10081 1317 10115
rect 1351 10112 1363 10115
rect 1504 10112 1532 10220
rect 2682 10208 2688 10220
rect 2740 10248 2746 10260
rect 3237 10251 3295 10257
rect 3237 10248 3249 10251
rect 2740 10220 3249 10248
rect 2740 10208 2746 10220
rect 3237 10217 3249 10220
rect 3283 10217 3295 10251
rect 3510 10248 3516 10260
rect 3237 10211 3295 10217
rect 3436 10220 3516 10248
rect 2866 10140 2872 10192
rect 2924 10180 2930 10192
rect 2924 10152 3188 10180
rect 2924 10140 2930 10152
rect 1351 10084 1532 10112
rect 1581 10115 1639 10121
rect 1351 10081 1363 10084
rect 1305 10075 1363 10081
rect 1581 10081 1593 10115
rect 1627 10112 1639 10115
rect 2406 10112 2412 10124
rect 1627 10084 2412 10112
rect 1627 10081 1639 10084
rect 1581 10075 1639 10081
rect 2406 10072 2412 10084
rect 2464 10072 2470 10124
rect 2774 10072 2780 10124
rect 2832 10121 2838 10124
rect 3160 10121 3188 10152
rect 3436 10124 3464 10220
rect 3510 10208 3516 10220
rect 3568 10248 3574 10260
rect 3694 10248 3700 10260
rect 3568 10220 3700 10248
rect 3568 10208 3574 10220
rect 3694 10208 3700 10220
rect 3752 10248 3758 10260
rect 5169 10251 5227 10257
rect 3752 10220 5120 10248
rect 3752 10208 3758 10220
rect 4556 10183 4614 10189
rect 4556 10149 4568 10183
rect 4602 10180 4614 10183
rect 4982 10180 4988 10192
rect 4602 10152 4988 10180
rect 4602 10149 4614 10152
rect 4556 10143 4614 10149
rect 4982 10140 4988 10152
rect 5040 10140 5046 10192
rect 2832 10075 2844 10121
rect 3145 10115 3203 10121
rect 3145 10081 3157 10115
rect 3191 10081 3203 10115
rect 3145 10075 3203 10081
rect 3329 10115 3387 10121
rect 3329 10081 3341 10115
rect 3375 10112 3387 10115
rect 3418 10112 3424 10124
rect 3375 10084 3424 10112
rect 3375 10081 3387 10084
rect 3329 10075 3387 10081
rect 2832 10072 2838 10075
rect 3418 10072 3424 10084
rect 3476 10072 3482 10124
rect 4154 10072 4160 10124
rect 4212 10112 4218 10124
rect 5092 10121 5120 10220
rect 5169 10217 5181 10251
rect 5215 10248 5227 10251
rect 5350 10248 5356 10260
rect 5215 10220 5356 10248
rect 5215 10217 5227 10220
rect 5169 10211 5227 10217
rect 5350 10208 5356 10220
rect 5408 10208 5414 10260
rect 7558 10248 7564 10260
rect 6840 10220 7564 10248
rect 6730 10180 6736 10192
rect 5644 10152 6736 10180
rect 4893 10115 4951 10121
rect 4893 10112 4905 10115
rect 4212 10084 4905 10112
rect 4212 10072 4218 10084
rect 4893 10081 4905 10084
rect 4939 10081 4951 10115
rect 4893 10075 4951 10081
rect 5077 10115 5135 10121
rect 5077 10081 5089 10115
rect 5123 10081 5135 10115
rect 5077 10075 5135 10081
rect 5353 10115 5411 10121
rect 5353 10081 5365 10115
rect 5399 10081 5411 10115
rect 5353 10075 5411 10081
rect 3050 10004 3056 10056
rect 3108 10004 3114 10056
rect 4798 10004 4804 10056
rect 4856 10004 4862 10056
rect 4985 10047 5043 10053
rect 4985 10013 4997 10047
rect 5031 10044 5043 10047
rect 5368 10044 5396 10075
rect 5534 10072 5540 10124
rect 5592 10072 5598 10124
rect 5644 10121 5672 10152
rect 6730 10140 6736 10152
rect 6788 10140 6794 10192
rect 5629 10115 5687 10121
rect 5629 10081 5641 10115
rect 5675 10081 5687 10115
rect 5629 10075 5687 10081
rect 5997 10115 6055 10121
rect 5997 10081 6009 10115
rect 6043 10112 6055 10115
rect 6840 10112 6868 10220
rect 7558 10208 7564 10220
rect 7616 10208 7622 10260
rect 8110 10208 8116 10260
rect 8168 10248 8174 10260
rect 8573 10251 8631 10257
rect 8573 10248 8585 10251
rect 8168 10220 8585 10248
rect 8168 10208 8174 10220
rect 8573 10217 8585 10220
rect 8619 10217 8631 10251
rect 8573 10211 8631 10217
rect 9490 10208 9496 10260
rect 9548 10208 9554 10260
rect 9582 10208 9588 10260
rect 9640 10248 9646 10260
rect 9640 10220 10824 10248
rect 9640 10208 9646 10220
rect 9674 10180 9680 10192
rect 7116 10152 9680 10180
rect 6043 10084 6868 10112
rect 6043 10081 6055 10084
rect 5997 10075 6055 10081
rect 7006 10072 7012 10124
rect 7064 10072 7070 10124
rect 7116 10121 7144 10152
rect 9674 10140 9680 10152
rect 9732 10140 9738 10192
rect 7101 10115 7159 10121
rect 7101 10081 7113 10115
rect 7147 10081 7159 10115
rect 7101 10075 7159 10081
rect 7368 10115 7426 10121
rect 7368 10081 7380 10115
rect 7414 10112 7426 10115
rect 7650 10112 7656 10124
rect 7414 10084 7656 10112
rect 7414 10081 7426 10084
rect 7368 10075 7426 10081
rect 7650 10072 7656 10084
rect 7708 10072 7714 10124
rect 7834 10072 7840 10124
rect 7892 10112 7898 10124
rect 7892 10084 8156 10112
rect 7892 10072 7898 10084
rect 5031 10016 5396 10044
rect 6273 10047 6331 10053
rect 5031 10013 5043 10016
rect 4985 10007 5043 10013
rect 6273 10013 6285 10047
rect 6319 10044 6331 10047
rect 6365 10047 6423 10053
rect 6365 10044 6377 10047
rect 6319 10016 6377 10044
rect 6319 10013 6331 10016
rect 6273 10007 6331 10013
rect 6365 10013 6377 10016
rect 6411 10013 6423 10047
rect 8128 10044 8156 10084
rect 8202 10072 8208 10124
rect 8260 10112 8266 10124
rect 10796 10121 10824 10220
rect 9125 10115 9183 10121
rect 9125 10112 9137 10115
rect 8260 10084 9137 10112
rect 8260 10072 8266 10084
rect 9125 10081 9137 10084
rect 9171 10081 9183 10115
rect 9125 10075 9183 10081
rect 9309 10115 9367 10121
rect 9309 10081 9321 10115
rect 9355 10081 9367 10115
rect 10597 10115 10655 10121
rect 10597 10112 10609 10115
rect 9309 10075 9367 10081
rect 10244 10084 10609 10112
rect 9324 10044 9352 10075
rect 10244 10053 10272 10084
rect 10597 10081 10609 10084
rect 10643 10081 10655 10115
rect 10597 10075 10655 10081
rect 10781 10115 10839 10121
rect 10781 10081 10793 10115
rect 10827 10081 10839 10115
rect 10781 10075 10839 10081
rect 8128 10016 9352 10044
rect 10229 10047 10287 10053
rect 6365 10007 6423 10013
rect 10229 10013 10241 10047
rect 10275 10013 10287 10047
rect 10229 10007 10287 10013
rect 1670 9936 1676 9988
rect 1728 9936 1734 9988
rect 6181 9979 6239 9985
rect 6181 9945 6193 9979
rect 6227 9976 6239 9979
rect 7098 9976 7104 9988
rect 6227 9948 7104 9976
rect 6227 9945 6239 9948
rect 6181 9939 6239 9945
rect 7098 9936 7104 9948
rect 7156 9936 7162 9988
rect 8294 9936 8300 9988
rect 8352 9976 8358 9988
rect 10244 9976 10272 10007
rect 10502 10004 10508 10056
rect 10560 10004 10566 10056
rect 8352 9948 10272 9976
rect 8352 9936 8358 9948
rect 1210 9868 1216 9920
rect 1268 9868 1274 9920
rect 1578 9868 1584 9920
rect 1636 9868 1642 9920
rect 3421 9911 3479 9917
rect 3421 9877 3433 9911
rect 3467 9908 3479 9911
rect 3602 9908 3608 9920
rect 3467 9880 3608 9908
rect 3467 9877 3479 9880
rect 3421 9871 3479 9877
rect 3602 9868 3608 9880
rect 3660 9908 3666 9920
rect 3878 9908 3884 9920
rect 3660 9880 3884 9908
rect 3660 9868 3666 9880
rect 3878 9868 3884 9880
rect 3936 9868 3942 9920
rect 5810 9868 5816 9920
rect 5868 9868 5874 9920
rect 7006 9868 7012 9920
rect 7064 9908 7070 9920
rect 7742 9908 7748 9920
rect 7064 9880 7748 9908
rect 7064 9868 7070 9880
rect 7742 9868 7748 9880
rect 7800 9868 7806 9920
rect 8018 9868 8024 9920
rect 8076 9908 8082 9920
rect 8481 9911 8539 9917
rect 8481 9908 8493 9911
rect 8076 9880 8493 9908
rect 8076 9868 8082 9880
rect 8481 9877 8493 9880
rect 8527 9877 8539 9911
rect 8481 9871 8539 9877
rect 9766 9868 9772 9920
rect 9824 9908 9830 9920
rect 10597 9911 10655 9917
rect 10597 9908 10609 9911
rect 9824 9880 10609 9908
rect 9824 9868 9830 9880
rect 10597 9877 10609 9880
rect 10643 9877 10655 9911
rect 10597 9871 10655 9877
rect 552 9818 11408 9840
rect 552 9766 1755 9818
rect 1807 9766 1819 9818
rect 1871 9766 1883 9818
rect 1935 9766 1947 9818
rect 1999 9766 2011 9818
rect 2063 9766 4469 9818
rect 4521 9766 4533 9818
rect 4585 9766 4597 9818
rect 4649 9766 4661 9818
rect 4713 9766 4725 9818
rect 4777 9766 7183 9818
rect 7235 9766 7247 9818
rect 7299 9766 7311 9818
rect 7363 9766 7375 9818
rect 7427 9766 7439 9818
rect 7491 9766 9897 9818
rect 9949 9766 9961 9818
rect 10013 9766 10025 9818
rect 10077 9766 10089 9818
rect 10141 9766 10153 9818
rect 10205 9766 11408 9818
rect 552 9744 11408 9766
rect 1302 9664 1308 9716
rect 1360 9664 1366 9716
rect 5261 9707 5319 9713
rect 2976 9676 4384 9704
rect 1118 9596 1124 9648
rect 1176 9596 1182 9648
rect 2869 9639 2927 9645
rect 2869 9605 2881 9639
rect 2915 9636 2927 9639
rect 2976 9636 3004 9676
rect 2915 9608 3004 9636
rect 2915 9605 2927 9608
rect 2869 9599 2927 9605
rect 3050 9596 3056 9648
rect 3108 9596 3114 9648
rect 4356 9636 4384 9676
rect 5261 9673 5273 9707
rect 5307 9704 5319 9707
rect 5307 9676 6592 9704
rect 5307 9673 5319 9676
rect 5261 9667 5319 9673
rect 4890 9636 4896 9648
rect 4356 9608 4896 9636
rect 4890 9596 4896 9608
rect 4948 9596 4954 9648
rect 4985 9639 5043 9645
rect 4985 9605 4997 9639
rect 5031 9636 5043 9639
rect 5442 9636 5448 9648
rect 5031 9608 5448 9636
rect 5031 9605 5043 9608
rect 4985 9599 5043 9605
rect 5442 9596 5448 9608
rect 5500 9596 5506 9648
rect 6564 9636 6592 9676
rect 7006 9664 7012 9716
rect 7064 9664 7070 9716
rect 7929 9707 7987 9713
rect 7929 9673 7941 9707
rect 7975 9704 7987 9707
rect 8202 9704 8208 9716
rect 7975 9676 8208 9704
rect 7975 9673 7987 9676
rect 7929 9667 7987 9673
rect 8202 9664 8208 9676
rect 8260 9664 8266 9716
rect 8849 9707 8907 9713
rect 8849 9673 8861 9707
rect 8895 9704 8907 9707
rect 8938 9704 8944 9716
rect 8895 9676 8944 9704
rect 8895 9673 8907 9676
rect 8849 9667 8907 9673
rect 8938 9664 8944 9676
rect 8996 9664 9002 9716
rect 7282 9636 7288 9648
rect 6564 9608 7288 9636
rect 7282 9596 7288 9608
rect 7340 9596 7346 9648
rect 7653 9639 7711 9645
rect 7653 9605 7665 9639
rect 7699 9636 7711 9639
rect 8294 9636 8300 9648
rect 7699 9608 7788 9636
rect 7699 9605 7711 9608
rect 7653 9599 7711 9605
rect 2685 9571 2743 9577
rect 2685 9537 2697 9571
rect 2731 9568 2743 9571
rect 3068 9568 3096 9596
rect 7760 9580 7788 9608
rect 7852 9608 8300 9636
rect 4798 9568 4804 9580
rect 2731 9540 3464 9568
rect 2731 9537 2743 9540
rect 2685 9531 2743 9537
rect 1213 9503 1271 9509
rect 1213 9469 1225 9503
rect 1259 9469 1271 9503
rect 1213 9463 1271 9469
rect 1228 9364 1256 9463
rect 1578 9460 1584 9512
rect 1636 9500 1642 9512
rect 2418 9503 2476 9509
rect 2418 9500 2430 9503
rect 1636 9472 2430 9500
rect 1636 9460 1642 9472
rect 2418 9469 2430 9472
rect 2464 9469 2476 9503
rect 2418 9463 2476 9469
rect 3050 9460 3056 9512
rect 3108 9460 3114 9512
rect 3436 9509 3464 9540
rect 4448 9540 4804 9568
rect 3421 9503 3479 9509
rect 3421 9469 3433 9503
rect 3467 9500 3479 9503
rect 3510 9500 3516 9512
rect 3467 9472 3516 9500
rect 3467 9469 3479 9472
rect 3421 9463 3479 9469
rect 3510 9460 3516 9472
rect 3568 9500 3574 9512
rect 4448 9500 4476 9540
rect 4798 9528 4804 9540
rect 4856 9568 4862 9580
rect 5629 9571 5687 9577
rect 5629 9568 5641 9571
rect 4856 9540 5641 9568
rect 4856 9528 4862 9540
rect 5629 9537 5641 9540
rect 5675 9537 5687 9571
rect 5629 9531 5687 9537
rect 7742 9528 7748 9580
rect 7800 9528 7806 9580
rect 3568 9472 4476 9500
rect 5169 9503 5227 9509
rect 3568 9460 3574 9472
rect 5169 9469 5181 9503
rect 5215 9500 5227 9503
rect 5442 9500 5448 9512
rect 5215 9472 5448 9500
rect 5215 9469 5227 9472
rect 5169 9463 5227 9469
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 5537 9503 5595 9509
rect 5537 9469 5549 9503
rect 5583 9500 5595 9503
rect 7377 9503 7435 9509
rect 7377 9500 7389 9503
rect 5583 9472 7389 9500
rect 5583 9469 5595 9472
rect 5537 9463 5595 9469
rect 7377 9469 7389 9472
rect 7423 9500 7435 9503
rect 7576 9500 7696 9502
rect 7852 9500 7880 9608
rect 8294 9596 8300 9608
rect 8352 9636 8358 9648
rect 8481 9639 8539 9645
rect 8481 9636 8493 9639
rect 8352 9608 8493 9636
rect 8352 9596 8358 9608
rect 8481 9605 8493 9608
rect 8527 9605 8539 9639
rect 8481 9599 8539 9605
rect 10321 9639 10379 9645
rect 10321 9605 10333 9639
rect 10367 9636 10379 9639
rect 10594 9636 10600 9648
rect 10367 9608 10600 9636
rect 10367 9605 10379 9608
rect 10321 9599 10379 9605
rect 10594 9596 10600 9608
rect 10652 9636 10658 9648
rect 10652 9608 11008 9636
rect 10652 9596 10658 9608
rect 10980 9577 11008 9608
rect 10965 9571 11023 9577
rect 10965 9537 10977 9571
rect 11011 9537 11023 9571
rect 10965 9531 11023 9537
rect 8389 9503 8447 9509
rect 8389 9500 8401 9503
rect 7423 9474 7880 9500
rect 7423 9472 7604 9474
rect 7668 9472 7880 9474
rect 8036 9472 8401 9500
rect 7423 9469 7435 9472
rect 7377 9463 7435 9469
rect 3326 9392 3332 9444
rect 3384 9432 3390 9444
rect 3666 9435 3724 9441
rect 3666 9432 3678 9435
rect 3384 9404 3678 9432
rect 3384 9392 3390 9404
rect 3666 9401 3678 9404
rect 3712 9401 3724 9435
rect 3666 9395 3724 9401
rect 4890 9392 4896 9444
rect 4948 9432 4954 9444
rect 5258 9432 5264 9444
rect 4948 9404 5264 9432
rect 4948 9392 4954 9404
rect 5258 9392 5264 9404
rect 5316 9392 5322 9444
rect 5902 9441 5908 9444
rect 5896 9395 5908 9441
rect 5902 9392 5908 9395
rect 5960 9392 5966 9444
rect 7469 9435 7527 9441
rect 7024 9404 7420 9432
rect 2590 9364 2596 9376
rect 1228 9336 2596 9364
rect 2590 9324 2596 9336
rect 2648 9324 2654 9376
rect 4062 9324 4068 9376
rect 4120 9364 4126 9376
rect 4801 9367 4859 9373
rect 4801 9364 4813 9367
rect 4120 9336 4813 9364
rect 4120 9324 4126 9336
rect 4801 9333 4813 9336
rect 4847 9333 4859 9367
rect 4801 9327 4859 9333
rect 5445 9367 5503 9373
rect 5445 9333 5457 9367
rect 5491 9364 5503 9367
rect 7024 9364 7052 9404
rect 5491 9336 7052 9364
rect 5491 9333 5503 9336
rect 5445 9327 5503 9333
rect 7098 9324 7104 9376
rect 7156 9324 7162 9376
rect 7282 9324 7288 9376
rect 7340 9324 7346 9376
rect 7392 9364 7420 9404
rect 7469 9401 7481 9435
rect 7515 9432 7527 9435
rect 7558 9432 7564 9444
rect 7515 9404 7564 9432
rect 7515 9401 7527 9404
rect 7469 9395 7527 9401
rect 7558 9392 7564 9404
rect 7616 9392 7622 9444
rect 8036 9432 8064 9472
rect 8389 9469 8401 9472
rect 8435 9469 8447 9503
rect 8389 9463 8447 9469
rect 7668 9404 8064 9432
rect 7668 9364 7696 9404
rect 8110 9392 8116 9444
rect 8168 9392 8174 9444
rect 7392 9336 7696 9364
rect 7742 9324 7748 9376
rect 7800 9324 7806 9376
rect 7913 9367 7971 9373
rect 7913 9333 7925 9367
rect 7959 9364 7971 9367
rect 8018 9364 8024 9376
rect 7959 9336 8024 9364
rect 7959 9333 7971 9336
rect 7913 9327 7971 9333
rect 8018 9324 8024 9336
rect 8076 9324 8082 9376
rect 8404 9364 8432 9463
rect 8662 9460 8668 9512
rect 8720 9460 8726 9512
rect 8941 9503 8999 9509
rect 8941 9469 8953 9503
rect 8987 9500 8999 9503
rect 9674 9500 9680 9512
rect 8987 9472 9680 9500
rect 8987 9469 8999 9472
rect 8941 9463 8999 9469
rect 9674 9460 9680 9472
rect 9732 9500 9738 9512
rect 10318 9500 10324 9512
rect 9732 9472 10324 9500
rect 9732 9460 9738 9472
rect 10318 9460 10324 9472
rect 10376 9460 10382 9512
rect 9030 9392 9036 9444
rect 9088 9432 9094 9444
rect 9186 9435 9244 9441
rect 9186 9432 9198 9435
rect 9088 9404 9198 9432
rect 9088 9392 9094 9404
rect 9186 9401 9198 9404
rect 9232 9401 9244 9435
rect 9186 9395 9244 9401
rect 10226 9364 10232 9376
rect 8404 9336 10232 9364
rect 10226 9324 10232 9336
rect 10284 9324 10290 9376
rect 10410 9324 10416 9376
rect 10468 9324 10474 9376
rect 552 9274 11568 9296
rect 552 9222 3112 9274
rect 3164 9222 3176 9274
rect 3228 9222 3240 9274
rect 3292 9222 3304 9274
rect 3356 9222 3368 9274
rect 3420 9222 5826 9274
rect 5878 9222 5890 9274
rect 5942 9222 5954 9274
rect 6006 9222 6018 9274
rect 6070 9222 6082 9274
rect 6134 9222 8540 9274
rect 8592 9222 8604 9274
rect 8656 9222 8668 9274
rect 8720 9222 8732 9274
rect 8784 9222 8796 9274
rect 8848 9222 11254 9274
rect 11306 9222 11318 9274
rect 11370 9222 11382 9274
rect 11434 9222 11446 9274
rect 11498 9222 11510 9274
rect 11562 9222 11568 9274
rect 552 9200 11568 9222
rect 2406 9120 2412 9172
rect 2464 9120 2470 9172
rect 2866 9160 2872 9172
rect 2746 9132 2872 9160
rect 2593 9027 2651 9033
rect 2593 8993 2605 9027
rect 2639 9024 2651 9027
rect 2746 9024 2774 9132
rect 2866 9120 2872 9132
rect 2924 9160 2930 9172
rect 3237 9163 3295 9169
rect 3237 9160 3249 9163
rect 2924 9132 3249 9160
rect 2924 9120 2930 9132
rect 3237 9129 3249 9132
rect 3283 9129 3295 9163
rect 3237 9123 3295 9129
rect 3405 9163 3463 9169
rect 3405 9129 3417 9163
rect 3451 9160 3463 9163
rect 3786 9160 3792 9172
rect 3451 9132 3792 9160
rect 3451 9129 3463 9132
rect 3405 9123 3463 9129
rect 3786 9120 3792 9132
rect 3844 9120 3850 9172
rect 5718 9120 5724 9172
rect 5776 9160 5782 9172
rect 5813 9163 5871 9169
rect 5813 9160 5825 9163
rect 5776 9132 5825 9160
rect 5776 9120 5782 9132
rect 5813 9129 5825 9132
rect 5859 9129 5871 9163
rect 5813 9123 5871 9129
rect 6549 9163 6607 9169
rect 6549 9129 6561 9163
rect 6595 9129 6607 9163
rect 6549 9123 6607 9129
rect 8021 9163 8079 9169
rect 8021 9129 8033 9163
rect 8067 9160 8079 9163
rect 9030 9160 9036 9172
rect 8067 9132 9036 9160
rect 8067 9129 8079 9132
rect 8021 9123 8079 9129
rect 3605 9095 3663 9101
rect 3605 9061 3617 9095
rect 3651 9092 3663 9095
rect 3970 9092 3976 9104
rect 3651 9064 3976 9092
rect 3651 9061 3663 9064
rect 3605 9055 3663 9061
rect 3970 9052 3976 9064
rect 4028 9052 4034 9104
rect 5445 9095 5503 9101
rect 5445 9061 5457 9095
rect 5491 9092 5503 9095
rect 6564 9092 6592 9123
rect 9030 9120 9036 9132
rect 9088 9120 9094 9172
rect 8573 9095 8631 9101
rect 8573 9092 8585 9095
rect 5491 9064 8585 9092
rect 5491 9061 5503 9064
rect 5445 9055 5503 9061
rect 8573 9061 8585 9064
rect 8619 9061 8631 9095
rect 8573 9055 8631 9061
rect 10318 9052 10324 9104
rect 10376 9092 10382 9104
rect 11054 9092 11060 9104
rect 10376 9064 11060 9092
rect 10376 9052 10382 9064
rect 11054 9052 11060 9064
rect 11112 9052 11118 9104
rect 2639 8996 2774 9024
rect 2869 9027 2927 9033
rect 2639 8993 2651 8996
rect 2593 8987 2651 8993
rect 2869 8993 2881 9027
rect 2915 9024 2927 9027
rect 4154 9024 4160 9036
rect 2915 8996 4160 9024
rect 2915 8993 2927 8996
rect 2869 8987 2927 8993
rect 4154 8984 4160 8996
rect 4212 8984 4218 9036
rect 5997 9027 6055 9033
rect 5997 8993 6009 9027
rect 6043 9024 6055 9027
rect 6362 9024 6368 9036
rect 6043 8996 6368 9024
rect 6043 8993 6055 8996
rect 5997 8987 6055 8993
rect 6362 8984 6368 8996
rect 6420 8984 6426 9036
rect 7834 8984 7840 9036
rect 7892 8984 7898 9036
rect 8205 9027 8263 9033
rect 8205 8993 8217 9027
rect 8251 8993 8263 9027
rect 8205 8987 8263 8993
rect 8481 9027 8539 9033
rect 8481 8993 8493 9027
rect 8527 9024 8539 9027
rect 10410 9024 10416 9036
rect 8527 8996 10416 9024
rect 8527 8993 8539 8996
rect 8481 8987 8539 8993
rect 2685 8959 2743 8965
rect 2685 8956 2697 8959
rect 2516 8928 2697 8956
rect 2516 8820 2544 8928
rect 2685 8925 2697 8928
rect 2731 8925 2743 8959
rect 2685 8919 2743 8925
rect 2777 8959 2835 8965
rect 2777 8925 2789 8959
rect 2823 8925 2835 8959
rect 2777 8919 2835 8925
rect 2590 8848 2596 8900
rect 2648 8888 2654 8900
rect 2792 8888 2820 8919
rect 3694 8916 3700 8968
rect 3752 8916 3758 8968
rect 5442 8916 5448 8968
rect 5500 8956 5506 8968
rect 7926 8956 7932 8968
rect 5500 8928 7932 8956
rect 5500 8916 5506 8928
rect 7926 8916 7932 8928
rect 7984 8916 7990 8968
rect 8220 8956 8248 8987
rect 10410 8984 10416 8996
rect 10468 8984 10474 9036
rect 10597 9027 10655 9033
rect 10597 8993 10609 9027
rect 10643 8993 10655 9027
rect 10597 8987 10655 8993
rect 9766 8956 9772 8968
rect 8220 8928 9772 8956
rect 9766 8916 9772 8928
rect 9824 8916 9830 8968
rect 10226 8916 10232 8968
rect 10284 8956 10290 8968
rect 10612 8956 10640 8987
rect 10284 8928 10640 8956
rect 10284 8916 10290 8928
rect 10778 8916 10784 8968
rect 10836 8916 10842 8968
rect 2648 8860 2820 8888
rect 2648 8848 2654 8860
rect 3326 8820 3332 8832
rect 2516 8792 3332 8820
rect 3326 8780 3332 8792
rect 3384 8780 3390 8832
rect 3421 8823 3479 8829
rect 3421 8789 3433 8823
rect 3467 8820 3479 8823
rect 4062 8820 4068 8832
rect 3467 8792 4068 8820
rect 3467 8789 3479 8792
rect 3421 8783 3479 8789
rect 4062 8780 4068 8792
rect 4120 8780 4126 8832
rect 7650 8780 7656 8832
rect 7708 8820 7714 8832
rect 8110 8820 8116 8832
rect 7708 8792 8116 8820
rect 7708 8780 7714 8792
rect 8110 8780 8116 8792
rect 8168 8780 8174 8832
rect 8294 8780 8300 8832
rect 8352 8820 8358 8832
rect 8389 8823 8447 8829
rect 8389 8820 8401 8823
rect 8352 8792 8401 8820
rect 8352 8780 8358 8792
rect 8389 8789 8401 8792
rect 8435 8789 8447 8823
rect 8389 8783 8447 8789
rect 10410 8780 10416 8832
rect 10468 8780 10474 8832
rect 552 8730 11408 8752
rect 552 8678 1755 8730
rect 1807 8678 1819 8730
rect 1871 8678 1883 8730
rect 1935 8678 1947 8730
rect 1999 8678 2011 8730
rect 2063 8678 4469 8730
rect 4521 8678 4533 8730
rect 4585 8678 4597 8730
rect 4649 8678 4661 8730
rect 4713 8678 4725 8730
rect 4777 8678 7183 8730
rect 7235 8678 7247 8730
rect 7299 8678 7311 8730
rect 7363 8678 7375 8730
rect 7427 8678 7439 8730
rect 7491 8678 9897 8730
rect 9949 8678 9961 8730
rect 10013 8678 10025 8730
rect 10077 8678 10089 8730
rect 10141 8678 10153 8730
rect 10205 8678 11408 8730
rect 552 8656 11408 8678
rect 2774 8576 2780 8628
rect 2832 8616 2838 8628
rect 2869 8619 2927 8625
rect 2869 8616 2881 8619
rect 2832 8588 2881 8616
rect 2832 8576 2838 8588
rect 2869 8585 2881 8588
rect 2915 8585 2927 8619
rect 4249 8619 4307 8625
rect 4249 8616 4261 8619
rect 2869 8579 2927 8585
rect 3344 8588 4261 8616
rect 2958 8372 2964 8424
rect 3016 8412 3022 8424
rect 3053 8415 3111 8421
rect 3053 8412 3065 8415
rect 3016 8384 3065 8412
rect 3016 8372 3022 8384
rect 3053 8381 3065 8384
rect 3099 8381 3111 8415
rect 3053 8375 3111 8381
rect 3237 8415 3295 8421
rect 3237 8381 3249 8415
rect 3283 8412 3295 8415
rect 3344 8412 3372 8588
rect 4249 8585 4261 8588
rect 4295 8585 4307 8619
rect 4249 8579 4307 8585
rect 7006 8576 7012 8628
rect 7064 8616 7070 8628
rect 7469 8619 7527 8625
rect 7469 8616 7481 8619
rect 7064 8588 7481 8616
rect 7064 8576 7070 8588
rect 7469 8585 7481 8588
rect 7515 8585 7527 8619
rect 7469 8579 7527 8585
rect 3421 8551 3479 8557
rect 3421 8517 3433 8551
rect 3467 8548 3479 8551
rect 3510 8548 3516 8560
rect 3467 8520 3516 8548
rect 3467 8517 3479 8520
rect 3421 8511 3479 8517
rect 3510 8508 3516 8520
rect 3568 8508 3574 8560
rect 4062 8548 4068 8560
rect 3712 8520 4068 8548
rect 3712 8480 3740 8520
rect 4062 8508 4068 8520
rect 4120 8508 4126 8560
rect 4157 8551 4215 8557
rect 4157 8517 4169 8551
rect 4203 8548 4215 8551
rect 5166 8548 5172 8560
rect 4203 8520 5172 8548
rect 4203 8517 4215 8520
rect 4157 8511 4215 8517
rect 5166 8508 5172 8520
rect 5224 8508 5230 8560
rect 6365 8551 6423 8557
rect 6365 8548 6377 8551
rect 5736 8520 6377 8548
rect 4706 8480 4712 8492
rect 3528 8452 3740 8480
rect 3804 8452 4712 8480
rect 3528 8421 3556 8452
rect 3283 8384 3372 8412
rect 3421 8415 3479 8421
rect 3283 8381 3295 8384
rect 3237 8375 3295 8381
rect 3421 8381 3433 8415
rect 3467 8412 3479 8415
rect 3513 8415 3571 8421
rect 3513 8412 3525 8415
rect 3467 8384 3525 8412
rect 3467 8381 3479 8384
rect 3421 8375 3479 8381
rect 3513 8381 3525 8384
rect 3559 8381 3571 8415
rect 3513 8375 3571 8381
rect 2958 8236 2964 8288
rect 3016 8276 3022 8288
rect 3252 8276 3280 8375
rect 3602 8372 3608 8424
rect 3660 8412 3666 8424
rect 3804 8421 3832 8452
rect 4706 8440 4712 8452
rect 4764 8440 4770 8492
rect 5629 8483 5687 8489
rect 5629 8480 5641 8483
rect 4816 8452 5641 8480
rect 3697 8415 3755 8421
rect 3697 8412 3709 8415
rect 3660 8384 3709 8412
rect 3660 8372 3666 8384
rect 3697 8381 3709 8384
rect 3743 8381 3755 8415
rect 3697 8375 3755 8381
rect 3789 8415 3847 8421
rect 3789 8381 3801 8415
rect 3835 8381 3847 8415
rect 3789 8375 3847 8381
rect 3881 8415 3939 8421
rect 3881 8381 3893 8415
rect 3927 8381 3939 8415
rect 3881 8375 3939 8381
rect 3326 8304 3332 8356
rect 3384 8344 3390 8356
rect 3896 8344 3924 8375
rect 3970 8372 3976 8424
rect 4028 8372 4034 8424
rect 4816 8412 4844 8452
rect 5629 8449 5641 8452
rect 5675 8449 5687 8483
rect 5629 8443 5687 8449
rect 5736 8424 5764 8520
rect 6365 8517 6377 8520
rect 6411 8548 6423 8551
rect 7484 8548 7512 8579
rect 7742 8576 7748 8628
rect 7800 8616 7806 8628
rect 8757 8619 8815 8625
rect 8757 8616 8769 8619
rect 7800 8588 8769 8616
rect 7800 8576 7806 8588
rect 8757 8585 8769 8588
rect 8803 8585 8815 8619
rect 8757 8579 8815 8585
rect 8113 8551 8171 8557
rect 8113 8548 8125 8551
rect 6411 8520 7328 8548
rect 7484 8520 8125 8548
rect 6411 8517 6423 8520
rect 6365 8511 6423 8517
rect 7098 8480 7104 8492
rect 5828 8452 7104 8480
rect 4080 8384 4844 8412
rect 4893 8415 4951 8421
rect 4080 8344 4108 8384
rect 4893 8381 4905 8415
rect 4939 8381 4951 8415
rect 4893 8375 4951 8381
rect 5537 8415 5595 8421
rect 5537 8381 5549 8415
rect 5583 8412 5595 8415
rect 5718 8412 5724 8424
rect 5583 8384 5724 8412
rect 5583 8381 5595 8384
rect 5537 8375 5595 8381
rect 3384 8316 4108 8344
rect 3384 8304 3390 8316
rect 4154 8304 4160 8356
rect 4212 8344 4218 8356
rect 4798 8344 4804 8356
rect 4212 8316 4804 8344
rect 4212 8304 4218 8316
rect 4798 8304 4804 8316
rect 4856 8304 4862 8356
rect 4908 8344 4936 8375
rect 5718 8372 5724 8384
rect 5776 8372 5782 8424
rect 5828 8421 5856 8452
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 5813 8415 5871 8421
rect 5813 8381 5825 8415
rect 5859 8381 5871 8415
rect 5813 8375 5871 8381
rect 6181 8415 6239 8421
rect 6181 8381 6193 8415
rect 6227 8412 6239 8415
rect 6270 8412 6276 8424
rect 6227 8384 6276 8412
rect 6227 8381 6239 8384
rect 6181 8375 6239 8381
rect 6270 8372 6276 8384
rect 6328 8372 6334 8424
rect 6454 8372 6460 8424
rect 6512 8372 6518 8424
rect 6733 8415 6791 8421
rect 6733 8381 6745 8415
rect 6779 8381 6791 8415
rect 6733 8375 6791 8381
rect 4982 8344 4988 8356
rect 4908 8316 4988 8344
rect 4982 8304 4988 8316
rect 5040 8304 5046 8356
rect 5074 8304 5080 8356
rect 5132 8344 5138 8356
rect 5353 8347 5411 8353
rect 5353 8344 5365 8347
rect 5132 8316 5365 8344
rect 5132 8304 5138 8316
rect 5353 8313 5365 8316
rect 5399 8313 5411 8347
rect 5353 8307 5411 8313
rect 6549 8347 6607 8353
rect 6549 8313 6561 8347
rect 6595 8344 6607 8347
rect 6638 8344 6644 8356
rect 6595 8316 6644 8344
rect 6595 8313 6607 8316
rect 6549 8307 6607 8313
rect 6638 8304 6644 8316
rect 6696 8304 6702 8356
rect 6748 8344 6776 8375
rect 6822 8372 6828 8424
rect 6880 8372 6886 8424
rect 6914 8372 6920 8424
rect 6972 8372 6978 8424
rect 7190 8372 7196 8424
rect 7248 8372 7254 8424
rect 7300 8421 7328 8520
rect 8113 8517 8125 8520
rect 8159 8517 8171 8551
rect 8113 8511 8171 8517
rect 7285 8415 7343 8421
rect 7285 8381 7297 8415
rect 7331 8412 7343 8415
rect 7466 8412 7472 8424
rect 7331 8384 7472 8412
rect 7331 8381 7343 8384
rect 7285 8375 7343 8381
rect 7466 8372 7472 8384
rect 7524 8372 7530 8424
rect 7742 8372 7748 8424
rect 7800 8372 7806 8424
rect 7926 8372 7932 8424
rect 7984 8372 7990 8424
rect 8202 8372 8208 8424
rect 8260 8372 8266 8424
rect 8573 8415 8631 8421
rect 8573 8381 8585 8415
rect 8619 8381 8631 8415
rect 8573 8375 8631 8381
rect 7760 8344 7788 8372
rect 6748 8316 7788 8344
rect 8386 8304 8392 8356
rect 8444 8304 8450 8356
rect 3016 8248 3280 8276
rect 3016 8236 3022 8248
rect 3786 8236 3792 8288
rect 3844 8236 3850 8288
rect 5166 8236 5172 8288
rect 5224 8236 5230 8288
rect 5258 8236 5264 8288
rect 5316 8236 5322 8288
rect 5997 8279 6055 8285
rect 5997 8245 6009 8279
rect 6043 8276 6055 8279
rect 6178 8276 6184 8288
rect 6043 8248 6184 8276
rect 6043 8245 6055 8248
rect 5997 8239 6055 8245
rect 6178 8236 6184 8248
rect 6236 8236 6242 8288
rect 6822 8236 6828 8288
rect 6880 8276 6886 8288
rect 7745 8279 7803 8285
rect 7745 8276 7757 8279
rect 6880 8248 7757 8276
rect 6880 8236 6886 8248
rect 7745 8245 7757 8248
rect 7791 8245 7803 8279
rect 8588 8276 8616 8375
rect 8846 8372 8852 8424
rect 8904 8372 8910 8424
rect 8941 8415 8999 8421
rect 8941 8381 8953 8415
rect 8987 8412 8999 8415
rect 9674 8412 9680 8424
rect 8987 8384 9680 8412
rect 8987 8381 8999 8384
rect 8941 8375 8999 8381
rect 9674 8372 9680 8384
rect 9732 8412 9738 8424
rect 10318 8412 10324 8424
rect 9732 8384 10324 8412
rect 9732 8372 9738 8384
rect 10318 8372 10324 8384
rect 10376 8372 10382 8424
rect 10962 8372 10968 8424
rect 11020 8372 11026 8424
rect 9030 8304 9036 8356
rect 9088 8344 9094 8356
rect 9186 8347 9244 8353
rect 9186 8344 9198 8347
rect 9088 8316 9198 8344
rect 9088 8304 9094 8316
rect 9186 8313 9198 8316
rect 9232 8313 9244 8347
rect 9186 8307 9244 8313
rect 9490 8304 9496 8356
rect 9548 8344 9554 8356
rect 10413 8347 10471 8353
rect 10413 8344 10425 8347
rect 9548 8316 10425 8344
rect 9548 8304 9554 8316
rect 10413 8313 10425 8316
rect 10459 8313 10471 8347
rect 10413 8307 10471 8313
rect 9306 8276 9312 8288
rect 8588 8248 9312 8276
rect 7745 8239 7803 8245
rect 9306 8236 9312 8248
rect 9364 8236 9370 8288
rect 10321 8279 10379 8285
rect 10321 8245 10333 8279
rect 10367 8276 10379 8279
rect 10962 8276 10968 8288
rect 10367 8248 10968 8276
rect 10367 8245 10379 8248
rect 10321 8239 10379 8245
rect 10962 8236 10968 8248
rect 11020 8236 11026 8288
rect 552 8186 11568 8208
rect 552 8134 3112 8186
rect 3164 8134 3176 8186
rect 3228 8134 3240 8186
rect 3292 8134 3304 8186
rect 3356 8134 3368 8186
rect 3420 8134 5826 8186
rect 5878 8134 5890 8186
rect 5942 8134 5954 8186
rect 6006 8134 6018 8186
rect 6070 8134 6082 8186
rect 6134 8134 8540 8186
rect 8592 8134 8604 8186
rect 8656 8134 8668 8186
rect 8720 8134 8732 8186
rect 8784 8134 8796 8186
rect 8848 8134 11254 8186
rect 11306 8134 11318 8186
rect 11370 8134 11382 8186
rect 11434 8134 11446 8186
rect 11498 8134 11510 8186
rect 11562 8134 11568 8186
rect 552 8112 11568 8134
rect 4706 8032 4712 8084
rect 4764 8072 4770 8084
rect 4801 8075 4859 8081
rect 4801 8072 4813 8075
rect 4764 8044 4813 8072
rect 4764 8032 4770 8044
rect 4801 8041 4813 8044
rect 4847 8041 4859 8075
rect 4801 8035 4859 8041
rect 6454 8032 6460 8084
rect 6512 8072 6518 8084
rect 6733 8075 6791 8081
rect 6733 8072 6745 8075
rect 6512 8044 6745 8072
rect 6512 8032 6518 8044
rect 6733 8041 6745 8044
rect 6779 8041 6791 8075
rect 6733 8035 6791 8041
rect 6914 8032 6920 8084
rect 6972 8072 6978 8084
rect 7469 8075 7527 8081
rect 7469 8072 7481 8075
rect 6972 8044 7481 8072
rect 6972 8032 6978 8044
rect 7469 8041 7481 8044
rect 7515 8041 7527 8075
rect 7469 8035 7527 8041
rect 7558 8032 7564 8084
rect 7616 8072 7622 8084
rect 8110 8072 8116 8084
rect 7616 8044 8116 8072
rect 7616 8032 7622 8044
rect 8110 8032 8116 8044
rect 8168 8072 8174 8084
rect 8389 8075 8447 8081
rect 8389 8072 8401 8075
rect 8168 8044 8401 8072
rect 8168 8032 8174 8044
rect 8389 8041 8401 8044
rect 8435 8041 8447 8075
rect 8389 8035 8447 8041
rect 8938 8032 8944 8084
rect 8996 8032 9002 8084
rect 10229 8075 10287 8081
rect 10229 8041 10241 8075
rect 10275 8072 10287 8075
rect 10502 8072 10508 8084
rect 10275 8044 10508 8072
rect 10275 8041 10287 8044
rect 10229 8035 10287 8041
rect 10502 8032 10508 8044
rect 10560 8032 10566 8084
rect 10594 8032 10600 8084
rect 10652 8032 10658 8084
rect 3694 8004 3700 8016
rect 3160 7976 3700 8004
rect 2774 7896 2780 7948
rect 2832 7896 2838 7948
rect 2958 7896 2964 7948
rect 3016 7936 3022 7948
rect 3160 7945 3188 7976
rect 3694 7964 3700 7976
rect 3752 7964 3758 8016
rect 7650 7964 7656 8016
rect 7708 8004 7714 8016
rect 8018 8004 8024 8016
rect 7708 7976 8024 8004
rect 7708 7964 7714 7976
rect 8018 7964 8024 7976
rect 8076 8004 8082 8016
rect 8481 8007 8539 8013
rect 8481 8004 8493 8007
rect 8076 7976 8493 8004
rect 8076 7964 8082 7976
rect 8481 7973 8493 7976
rect 8527 7973 8539 8007
rect 8481 7967 8539 7973
rect 8956 7976 10088 8004
rect 8956 7948 8984 7976
rect 3418 7945 3424 7948
rect 3053 7939 3111 7945
rect 3053 7936 3065 7939
rect 3016 7908 3065 7936
rect 3016 7896 3022 7908
rect 3053 7905 3065 7908
rect 3099 7905 3111 7939
rect 3053 7899 3111 7905
rect 3145 7939 3203 7945
rect 3145 7905 3157 7939
rect 3191 7905 3203 7939
rect 3412 7936 3424 7945
rect 3379 7908 3424 7936
rect 3145 7899 3203 7905
rect 3412 7899 3424 7908
rect 3418 7896 3424 7899
rect 3476 7896 3482 7948
rect 5258 7896 5264 7948
rect 5316 7936 5322 7948
rect 6365 7939 6423 7945
rect 6365 7936 6377 7939
rect 5316 7908 6377 7936
rect 5316 7896 5322 7908
rect 6365 7905 6377 7908
rect 6411 7905 6423 7939
rect 6365 7899 6423 7905
rect 7558 7896 7564 7948
rect 7616 7936 7622 7948
rect 7745 7939 7803 7945
rect 7745 7936 7757 7939
rect 7616 7908 7757 7936
rect 7616 7896 7622 7908
rect 7745 7905 7757 7908
rect 7791 7905 7803 7939
rect 7745 7899 7803 7905
rect 7837 7939 7895 7945
rect 7837 7905 7849 7939
rect 7883 7936 7895 7939
rect 8113 7939 8171 7945
rect 8113 7936 8125 7939
rect 7883 7908 8125 7936
rect 7883 7905 7895 7908
rect 7837 7899 7895 7905
rect 8113 7905 8125 7908
rect 8159 7905 8171 7939
rect 8113 7899 8171 7905
rect 8297 7939 8355 7945
rect 8297 7905 8309 7939
rect 8343 7905 8355 7939
rect 8297 7899 8355 7905
rect 5442 7828 5448 7880
rect 5500 7828 5506 7880
rect 7190 7828 7196 7880
rect 7248 7868 7254 7880
rect 7377 7871 7435 7877
rect 7377 7868 7389 7871
rect 7248 7840 7389 7868
rect 7248 7828 7254 7840
rect 7377 7837 7389 7840
rect 7423 7837 7435 7871
rect 7377 7831 7435 7837
rect 7392 7800 7420 7831
rect 7466 7828 7472 7880
rect 7524 7868 7530 7880
rect 7653 7871 7711 7877
rect 7653 7868 7665 7871
rect 7524 7840 7665 7868
rect 7524 7828 7530 7840
rect 7653 7837 7665 7840
rect 7699 7837 7711 7871
rect 7852 7868 7880 7899
rect 7653 7831 7711 7837
rect 7760 7840 7880 7868
rect 7929 7871 7987 7877
rect 7760 7812 7788 7840
rect 7929 7837 7941 7871
rect 7975 7868 7987 7871
rect 8202 7868 8208 7880
rect 7975 7840 8208 7868
rect 7975 7837 7987 7840
rect 7929 7831 7987 7837
rect 8202 7828 8208 7840
rect 8260 7828 8266 7880
rect 8312 7868 8340 7899
rect 8938 7896 8944 7948
rect 8996 7896 9002 7948
rect 9398 7896 9404 7948
rect 9456 7936 9462 7948
rect 10060 7945 10088 7976
rect 10410 7964 10416 8016
rect 10468 7964 10474 8016
rect 9861 7939 9919 7945
rect 9861 7936 9873 7939
rect 9456 7908 9873 7936
rect 9456 7896 9462 7908
rect 9861 7905 9873 7908
rect 9907 7905 9919 7939
rect 9861 7899 9919 7905
rect 10045 7939 10103 7945
rect 10045 7905 10057 7939
rect 10091 7936 10103 7939
rect 10505 7939 10563 7945
rect 10505 7936 10517 7939
rect 10091 7908 10517 7936
rect 10091 7905 10103 7908
rect 10045 7899 10103 7905
rect 10505 7905 10517 7908
rect 10551 7905 10563 7939
rect 10505 7899 10563 7905
rect 9122 7868 9128 7880
rect 8312 7840 9128 7868
rect 9122 7828 9128 7840
rect 9180 7868 9186 7880
rect 9493 7871 9551 7877
rect 9493 7868 9505 7871
rect 9180 7840 9505 7868
rect 9180 7828 9186 7840
rect 9493 7837 9505 7840
rect 9539 7837 9551 7871
rect 9493 7831 9551 7837
rect 9766 7828 9772 7880
rect 9824 7868 9830 7880
rect 10137 7871 10195 7877
rect 10137 7868 10149 7871
rect 9824 7840 10149 7868
rect 9824 7828 9830 7840
rect 10137 7837 10149 7840
rect 10183 7837 10195 7871
rect 11146 7868 11152 7880
rect 10137 7831 10195 7837
rect 10244 7840 11152 7868
rect 7742 7800 7748 7812
rect 7392 7772 7748 7800
rect 7742 7760 7748 7772
rect 7800 7760 7806 7812
rect 10244 7800 10272 7840
rect 11146 7828 11152 7840
rect 11204 7828 11210 7880
rect 7944 7772 10272 7800
rect 10781 7803 10839 7809
rect 2590 7692 2596 7744
rect 2648 7692 2654 7744
rect 2958 7692 2964 7744
rect 3016 7692 3022 7744
rect 3326 7692 3332 7744
rect 3384 7732 3390 7744
rect 4525 7735 4583 7741
rect 4525 7732 4537 7735
rect 3384 7704 4537 7732
rect 3384 7692 3390 7704
rect 4525 7701 4537 7704
rect 4571 7732 4583 7735
rect 4982 7732 4988 7744
rect 4571 7704 4988 7732
rect 4571 7701 4583 7704
rect 4525 7695 4583 7701
rect 4982 7692 4988 7704
rect 5040 7732 5046 7744
rect 5350 7732 5356 7744
rect 5040 7704 5356 7732
rect 5040 7692 5046 7704
rect 5350 7692 5356 7704
rect 5408 7692 5414 7744
rect 5534 7692 5540 7744
rect 5592 7732 5598 7744
rect 5813 7735 5871 7741
rect 5813 7732 5825 7735
rect 5592 7704 5825 7732
rect 5592 7692 5598 7704
rect 5813 7701 5825 7704
rect 5859 7701 5871 7735
rect 5813 7695 5871 7701
rect 6362 7692 6368 7744
rect 6420 7732 6426 7744
rect 7944 7732 7972 7772
rect 10781 7769 10793 7803
rect 10827 7800 10839 7803
rect 10962 7800 10968 7812
rect 10827 7772 10968 7800
rect 10827 7769 10839 7772
rect 10781 7763 10839 7769
rect 10962 7760 10968 7772
rect 11020 7760 11026 7812
rect 6420 7704 7972 7732
rect 8665 7735 8723 7741
rect 6420 7692 6426 7704
rect 8665 7701 8677 7735
rect 8711 7732 8723 7735
rect 9214 7732 9220 7744
rect 8711 7704 9220 7732
rect 8711 7701 8723 7704
rect 8665 7695 8723 7701
rect 9214 7692 9220 7704
rect 9272 7692 9278 7744
rect 9582 7692 9588 7744
rect 9640 7732 9646 7744
rect 9677 7735 9735 7741
rect 9677 7732 9689 7735
rect 9640 7704 9689 7732
rect 9640 7692 9646 7704
rect 9677 7701 9689 7704
rect 9723 7701 9735 7735
rect 9677 7695 9735 7701
rect 552 7642 11408 7664
rect 552 7590 1755 7642
rect 1807 7590 1819 7642
rect 1871 7590 1883 7642
rect 1935 7590 1947 7642
rect 1999 7590 2011 7642
rect 2063 7590 4469 7642
rect 4521 7590 4533 7642
rect 4585 7590 4597 7642
rect 4649 7590 4661 7642
rect 4713 7590 4725 7642
rect 4777 7590 7183 7642
rect 7235 7590 7247 7642
rect 7299 7590 7311 7642
rect 7363 7590 7375 7642
rect 7427 7590 7439 7642
rect 7491 7590 9897 7642
rect 9949 7590 9961 7642
rect 10013 7590 10025 7642
rect 10077 7590 10089 7642
rect 10141 7590 10153 7642
rect 10205 7590 11408 7642
rect 552 7568 11408 7590
rect 2409 7531 2467 7537
rect 2409 7497 2421 7531
rect 2455 7528 2467 7531
rect 2958 7528 2964 7540
rect 2455 7500 2964 7528
rect 2455 7497 2467 7500
rect 2409 7491 2467 7497
rect 2958 7488 2964 7500
rect 3016 7488 3022 7540
rect 3421 7531 3479 7537
rect 3421 7497 3433 7531
rect 3467 7528 3479 7531
rect 3510 7528 3516 7540
rect 3467 7500 3516 7528
rect 3467 7497 3479 7500
rect 3421 7491 3479 7497
rect 1765 7395 1823 7401
rect 1765 7361 1777 7395
rect 1811 7392 1823 7395
rect 2590 7392 2596 7404
rect 1811 7364 2596 7392
rect 1811 7361 1823 7364
rect 1765 7355 1823 7361
rect 2590 7352 2596 7364
rect 2648 7352 2654 7404
rect 3053 7395 3111 7401
rect 3053 7361 3065 7395
rect 3099 7392 3111 7395
rect 3436 7392 3464 7491
rect 3510 7488 3516 7500
rect 3568 7528 3574 7540
rect 5166 7528 5172 7540
rect 3568 7500 5172 7528
rect 3568 7488 3574 7500
rect 5166 7488 5172 7500
rect 5224 7488 5230 7540
rect 5442 7488 5448 7540
rect 5500 7488 5506 7540
rect 7009 7531 7067 7537
rect 7009 7497 7021 7531
rect 7055 7528 7067 7531
rect 7098 7528 7104 7540
rect 7055 7500 7104 7528
rect 7055 7497 7067 7500
rect 7009 7491 7067 7497
rect 7098 7488 7104 7500
rect 7156 7488 7162 7540
rect 7377 7531 7435 7537
rect 7377 7497 7389 7531
rect 7423 7528 7435 7531
rect 7926 7528 7932 7540
rect 7423 7500 7932 7528
rect 7423 7497 7435 7500
rect 7377 7491 7435 7497
rect 7926 7488 7932 7500
rect 7984 7488 7990 7540
rect 8202 7488 8208 7540
rect 8260 7488 8266 7540
rect 9306 7488 9312 7540
rect 9364 7488 9370 7540
rect 3099 7364 3464 7392
rect 3099 7361 3111 7364
rect 3053 7355 3111 7361
rect 9214 7352 9220 7404
rect 9272 7352 9278 7404
rect 10229 7395 10287 7401
rect 10229 7361 10241 7395
rect 10275 7392 10287 7395
rect 10778 7392 10784 7404
rect 10275 7364 10784 7392
rect 10275 7361 10287 7364
rect 10229 7355 10287 7361
rect 10778 7352 10784 7364
rect 10836 7352 10842 7404
rect 3694 7284 3700 7336
rect 3752 7284 3758 7336
rect 3786 7284 3792 7336
rect 3844 7324 3850 7336
rect 3953 7327 4011 7333
rect 3953 7324 3965 7327
rect 3844 7296 3965 7324
rect 3844 7284 3850 7296
rect 3953 7293 3965 7296
rect 3999 7293 4011 7327
rect 3953 7287 4011 7293
rect 5166 7284 5172 7336
rect 5224 7284 5230 7336
rect 5258 7284 5264 7336
rect 5316 7284 5322 7336
rect 5445 7327 5503 7333
rect 5445 7293 5457 7327
rect 5491 7324 5503 7327
rect 5534 7324 5540 7336
rect 5491 7296 5540 7324
rect 5491 7293 5503 7296
rect 5445 7287 5503 7293
rect 5534 7284 5540 7296
rect 5592 7284 5598 7336
rect 5626 7284 5632 7336
rect 5684 7284 5690 7336
rect 5896 7327 5954 7333
rect 5896 7293 5908 7327
rect 5942 7324 5954 7327
rect 6178 7324 6184 7336
rect 5942 7296 6184 7324
rect 5942 7293 5954 7296
rect 5896 7287 5954 7293
rect 6178 7284 6184 7296
rect 6236 7284 6242 7336
rect 7098 7284 7104 7336
rect 7156 7284 7162 7336
rect 7653 7327 7711 7333
rect 7653 7293 7665 7327
rect 7699 7324 7711 7327
rect 7742 7324 7748 7336
rect 7699 7296 7748 7324
rect 7699 7293 7711 7296
rect 7653 7287 7711 7293
rect 7742 7284 7748 7296
rect 7800 7284 7806 7336
rect 8938 7284 8944 7336
rect 8996 7324 9002 7336
rect 9309 7327 9367 7333
rect 9309 7324 9321 7327
rect 8996 7296 9321 7324
rect 8996 7284 9002 7296
rect 9309 7293 9321 7296
rect 9355 7293 9367 7327
rect 9309 7287 9367 7293
rect 9493 7327 9551 7333
rect 9493 7293 9505 7327
rect 9539 7293 9551 7327
rect 9493 7287 9551 7293
rect 10413 7327 10471 7333
rect 10413 7293 10425 7327
rect 10459 7324 10471 7327
rect 10502 7324 10508 7336
rect 10459 7296 10508 7324
rect 10459 7293 10471 7296
rect 10413 7287 10471 7293
rect 2317 7259 2375 7265
rect 2317 7225 2329 7259
rect 2363 7256 2375 7259
rect 2498 7256 2504 7268
rect 2363 7228 2504 7256
rect 2363 7225 2375 7228
rect 2317 7219 2375 7225
rect 2498 7216 2504 7228
rect 2556 7216 2562 7268
rect 2958 7216 2964 7268
rect 3016 7256 3022 7268
rect 3237 7259 3295 7265
rect 3237 7256 3249 7259
rect 3016 7228 3249 7256
rect 3016 7216 3022 7228
rect 3237 7225 3249 7228
rect 3283 7256 3295 7259
rect 3326 7256 3332 7268
rect 3283 7228 3332 7256
rect 3283 7225 3295 7228
rect 3237 7219 3295 7225
rect 3326 7216 3332 7228
rect 3384 7216 3390 7268
rect 3453 7259 3511 7265
rect 3453 7225 3465 7259
rect 3499 7256 3511 7259
rect 5276 7256 5304 7284
rect 3499 7228 5304 7256
rect 3499 7225 3511 7228
rect 3453 7219 3511 7225
rect 3602 7148 3608 7200
rect 3660 7148 3666 7200
rect 5092 7197 5120 7228
rect 6730 7216 6736 7268
rect 6788 7256 6794 7268
rect 7377 7259 7435 7265
rect 7377 7256 7389 7259
rect 6788 7228 7389 7256
rect 6788 7216 6794 7228
rect 7377 7225 7389 7228
rect 7423 7256 7435 7259
rect 7926 7256 7932 7268
rect 7423 7228 7932 7256
rect 7423 7225 7435 7228
rect 7377 7219 7435 7225
rect 7926 7216 7932 7228
rect 7984 7216 7990 7268
rect 8202 7216 8208 7268
rect 8260 7256 8266 7268
rect 9508 7256 9536 7287
rect 10502 7284 10508 7296
rect 10560 7284 10566 7336
rect 8260 7228 9536 7256
rect 8260 7216 8266 7228
rect 5077 7191 5135 7197
rect 5077 7157 5089 7191
rect 5123 7157 5135 7191
rect 5077 7151 5135 7157
rect 5261 7191 5319 7197
rect 5261 7157 5273 7191
rect 5307 7188 5319 7191
rect 5350 7188 5356 7200
rect 5307 7160 5356 7188
rect 5307 7157 5319 7160
rect 5261 7151 5319 7157
rect 5350 7148 5356 7160
rect 5408 7148 5414 7200
rect 7193 7191 7251 7197
rect 7193 7157 7205 7191
rect 7239 7188 7251 7191
rect 8110 7188 8116 7200
rect 7239 7160 8116 7188
rect 7239 7157 7251 7160
rect 7193 7151 7251 7157
rect 8110 7148 8116 7160
rect 8168 7148 8174 7200
rect 9214 7148 9220 7200
rect 9272 7188 9278 7200
rect 9585 7191 9643 7197
rect 9585 7188 9597 7191
rect 9272 7160 9597 7188
rect 9272 7148 9278 7160
rect 9585 7157 9597 7160
rect 9631 7188 9643 7191
rect 9766 7188 9772 7200
rect 9631 7160 9772 7188
rect 9631 7157 9643 7160
rect 9585 7151 9643 7157
rect 9766 7148 9772 7160
rect 9824 7148 9830 7200
rect 10686 7148 10692 7200
rect 10744 7188 10750 7200
rect 10965 7191 11023 7197
rect 10965 7188 10977 7191
rect 10744 7160 10977 7188
rect 10744 7148 10750 7160
rect 10965 7157 10977 7160
rect 11011 7157 11023 7191
rect 10965 7151 11023 7157
rect 552 7098 11568 7120
rect 552 7046 3112 7098
rect 3164 7046 3176 7098
rect 3228 7046 3240 7098
rect 3292 7046 3304 7098
rect 3356 7046 3368 7098
rect 3420 7046 5826 7098
rect 5878 7046 5890 7098
rect 5942 7046 5954 7098
rect 6006 7046 6018 7098
rect 6070 7046 6082 7098
rect 6134 7046 8540 7098
rect 8592 7046 8604 7098
rect 8656 7046 8668 7098
rect 8720 7046 8732 7098
rect 8784 7046 8796 7098
rect 8848 7046 11254 7098
rect 11306 7046 11318 7098
rect 11370 7046 11382 7098
rect 11434 7046 11446 7098
rect 11498 7046 11510 7098
rect 11562 7046 11568 7098
rect 552 7024 11568 7046
rect 3510 6944 3516 6996
rect 3568 6984 3574 6996
rect 3605 6987 3663 6993
rect 3605 6984 3617 6987
rect 3568 6956 3617 6984
rect 3568 6944 3574 6956
rect 3605 6953 3617 6956
rect 3651 6953 3663 6987
rect 3605 6947 3663 6953
rect 9122 6944 9128 6996
rect 9180 6984 9186 6996
rect 9217 6987 9275 6993
rect 9217 6984 9229 6987
rect 9180 6956 9229 6984
rect 9180 6944 9186 6956
rect 9217 6953 9229 6956
rect 9263 6953 9275 6987
rect 9217 6947 9275 6953
rect 10689 6987 10747 6993
rect 10689 6953 10701 6987
rect 10735 6984 10747 6987
rect 10778 6984 10784 6996
rect 10735 6956 10784 6984
rect 10735 6953 10747 6956
rect 10689 6947 10747 6953
rect 10778 6944 10784 6956
rect 10836 6944 10842 6996
rect 5626 6916 5632 6928
rect 2240 6888 5632 6916
rect 2240 6857 2268 6888
rect 2498 6857 2504 6860
rect 2225 6851 2283 6857
rect 2225 6817 2237 6851
rect 2271 6817 2283 6851
rect 2225 6811 2283 6817
rect 2492 6811 2504 6857
rect 2556 6848 2562 6860
rect 3896 6848 3924 6888
rect 5626 6876 5632 6888
rect 5684 6876 5690 6928
rect 7098 6916 7104 6928
rect 6472 6888 7104 6916
rect 3970 6857 3976 6860
rect 2556 6820 2592 6848
rect 3804 6820 3924 6848
rect 2498 6808 2504 6811
rect 2556 6808 2562 6820
rect 3694 6740 3700 6792
rect 3752 6780 3758 6792
rect 3804 6780 3832 6820
rect 3964 6811 3976 6857
rect 3970 6808 3976 6811
rect 4028 6808 4034 6860
rect 4246 6808 4252 6860
rect 4304 6848 4310 6860
rect 5169 6851 5227 6857
rect 5169 6848 5181 6851
rect 4304 6820 5181 6848
rect 4304 6808 4310 6820
rect 5169 6817 5181 6820
rect 5215 6817 5227 6851
rect 5169 6811 5227 6817
rect 5353 6851 5411 6857
rect 5353 6817 5365 6851
rect 5399 6848 5411 6851
rect 5718 6848 5724 6860
rect 5399 6820 5724 6848
rect 5399 6817 5411 6820
rect 5353 6811 5411 6817
rect 3752 6752 3832 6780
rect 5184 6780 5212 6811
rect 5718 6808 5724 6820
rect 5776 6808 5782 6860
rect 6086 6808 6092 6860
rect 6144 6808 6150 6860
rect 6273 6851 6331 6857
rect 6273 6817 6285 6851
rect 6319 6848 6331 6851
rect 6472 6848 6500 6888
rect 7098 6876 7104 6888
rect 7156 6876 7162 6928
rect 6638 6857 6644 6860
rect 6632 6848 6644 6857
rect 6319 6820 6500 6848
rect 6599 6820 6644 6848
rect 6319 6817 6331 6820
rect 6273 6811 6331 6817
rect 6632 6811 6644 6820
rect 6638 6808 6644 6811
rect 6696 6808 6702 6860
rect 8104 6851 8162 6857
rect 8104 6817 8116 6851
rect 8150 6848 8162 6851
rect 8386 6848 8392 6860
rect 8150 6820 8392 6848
rect 8150 6817 8162 6820
rect 8104 6811 8162 6817
rect 8386 6808 8392 6820
rect 8444 6808 8450 6860
rect 9582 6857 9588 6860
rect 9576 6848 9588 6857
rect 9543 6820 9588 6848
rect 9576 6811 9588 6820
rect 9582 6808 9588 6811
rect 9640 6808 9646 6860
rect 6095 6780 6123 6808
rect 5184 6752 6123 6780
rect 6365 6783 6423 6789
rect 3752 6740 3758 6752
rect 6365 6749 6377 6783
rect 6411 6749 6423 6783
rect 6365 6743 6423 6749
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6749 7895 6783
rect 7837 6743 7895 6749
rect 9309 6783 9367 6789
rect 9309 6749 9321 6783
rect 9355 6749 9367 6783
rect 9309 6743 9367 6749
rect 5074 6672 5080 6724
rect 5132 6672 5138 6724
rect 6270 6672 6276 6724
rect 6328 6672 6334 6724
rect 5350 6604 5356 6656
rect 5408 6604 5414 6656
rect 6380 6644 6408 6743
rect 7852 6712 7880 6743
rect 9324 6712 9352 6743
rect 7300 6684 7880 6712
rect 7300 6644 7328 6684
rect 6380 6616 7328 6644
rect 7742 6604 7748 6656
rect 7800 6604 7806 6656
rect 7852 6644 7880 6684
rect 8772 6684 9352 6712
rect 8772 6644 8800 6684
rect 7852 6616 8800 6644
rect 9324 6644 9352 6684
rect 9674 6644 9680 6656
rect 9324 6616 9680 6644
rect 9674 6604 9680 6616
rect 9732 6604 9738 6656
rect 552 6554 11408 6576
rect 552 6502 1755 6554
rect 1807 6502 1819 6554
rect 1871 6502 1883 6554
rect 1935 6502 1947 6554
rect 1999 6502 2011 6554
rect 2063 6502 4469 6554
rect 4521 6502 4533 6554
rect 4585 6502 4597 6554
rect 4649 6502 4661 6554
rect 4713 6502 4725 6554
rect 4777 6502 7183 6554
rect 7235 6502 7247 6554
rect 7299 6502 7311 6554
rect 7363 6502 7375 6554
rect 7427 6502 7439 6554
rect 7491 6502 9897 6554
rect 9949 6502 9961 6554
rect 10013 6502 10025 6554
rect 10077 6502 10089 6554
rect 10141 6502 10153 6554
rect 10205 6502 11408 6554
rect 552 6480 11408 6502
rect 2774 6400 2780 6452
rect 2832 6440 2838 6452
rect 3697 6443 3755 6449
rect 3697 6440 3709 6443
rect 2832 6412 3709 6440
rect 2832 6400 2838 6412
rect 3697 6409 3709 6412
rect 3743 6409 3755 6443
rect 3697 6403 3755 6409
rect 3970 6400 3976 6452
rect 4028 6440 4034 6452
rect 4157 6443 4215 6449
rect 4157 6440 4169 6443
rect 4028 6412 4169 6440
rect 4028 6400 4034 6412
rect 4157 6409 4169 6412
rect 4203 6409 4215 6443
rect 4157 6403 4215 6409
rect 6086 6400 6092 6452
rect 6144 6440 6150 6452
rect 6144 6412 7328 6440
rect 6144 6400 6150 6412
rect 3602 6332 3608 6384
rect 3660 6372 3666 6384
rect 4525 6375 4583 6381
rect 4525 6372 4537 6375
rect 3660 6344 4537 6372
rect 3660 6332 3666 6344
rect 4525 6341 4537 6344
rect 4571 6341 4583 6375
rect 4525 6335 4583 6341
rect 7193 6375 7251 6381
rect 7193 6341 7205 6375
rect 7239 6341 7251 6375
rect 7300 6372 7328 6412
rect 8110 6400 8116 6452
rect 8168 6400 8174 6452
rect 8941 6443 8999 6449
rect 8941 6409 8953 6443
rect 8987 6440 8999 6443
rect 9030 6440 9036 6452
rect 8987 6412 9036 6440
rect 8987 6409 8999 6412
rect 8941 6403 8999 6409
rect 9030 6400 9036 6412
rect 9088 6400 9094 6452
rect 9493 6443 9551 6449
rect 9493 6409 9505 6443
rect 9539 6440 9551 6443
rect 9858 6440 9864 6452
rect 9539 6412 9864 6440
rect 9539 6409 9551 6412
rect 9493 6403 9551 6409
rect 9858 6400 9864 6412
rect 9916 6440 9922 6452
rect 10226 6440 10232 6452
rect 9916 6412 10232 6440
rect 9916 6400 9922 6412
rect 10226 6400 10232 6412
rect 10284 6400 10290 6452
rect 8202 6372 8208 6384
rect 7300 6344 8208 6372
rect 7193 6335 7251 6341
rect 5350 6304 5356 6316
rect 4356 6276 5356 6304
rect 3510 6196 3516 6248
rect 3568 6236 3574 6248
rect 4356 6245 4384 6276
rect 5350 6264 5356 6276
rect 5408 6264 5414 6316
rect 5626 6264 5632 6316
rect 5684 6304 5690 6316
rect 5813 6307 5871 6313
rect 5813 6304 5825 6307
rect 5684 6276 5825 6304
rect 5684 6264 5690 6276
rect 5813 6273 5825 6276
rect 5859 6273 5871 6307
rect 7208 6304 7236 6335
rect 8202 6332 8208 6344
rect 8260 6372 8266 6384
rect 8386 6372 8392 6384
rect 8260 6344 8392 6372
rect 8260 6332 8266 6344
rect 8386 6332 8392 6344
rect 8444 6372 8450 6384
rect 8665 6375 8723 6381
rect 8665 6372 8677 6375
rect 8444 6344 8677 6372
rect 8444 6332 8450 6344
rect 8665 6341 8677 6344
rect 8711 6341 8723 6375
rect 8665 6335 8723 6341
rect 7558 6304 7564 6316
rect 7208 6276 7564 6304
rect 5813 6267 5871 6273
rect 7558 6264 7564 6276
rect 7616 6264 7622 6316
rect 9401 6307 9459 6313
rect 9401 6273 9413 6307
rect 9447 6304 9459 6307
rect 9490 6304 9496 6316
rect 9447 6276 9496 6304
rect 9447 6273 9459 6276
rect 9401 6267 9459 6273
rect 9490 6264 9496 6276
rect 9548 6264 9554 6316
rect 3973 6239 4031 6245
rect 3973 6236 3985 6239
rect 3568 6208 3985 6236
rect 3568 6196 3574 6208
rect 3973 6205 3985 6208
rect 4019 6205 4031 6239
rect 3973 6199 4031 6205
rect 4341 6239 4399 6245
rect 4341 6205 4353 6239
rect 4387 6205 4399 6239
rect 4341 6199 4399 6205
rect 4617 6239 4675 6245
rect 4617 6205 4629 6239
rect 4663 6236 4675 6239
rect 4893 6239 4951 6245
rect 4893 6236 4905 6239
rect 4663 6208 4905 6236
rect 4663 6205 4675 6208
rect 4617 6199 4675 6205
rect 4893 6205 4905 6208
rect 4939 6205 4951 6239
rect 4893 6199 4951 6205
rect 5074 6196 5080 6248
rect 5132 6236 5138 6248
rect 5445 6239 5503 6245
rect 5445 6236 5457 6239
rect 5132 6208 5457 6236
rect 5132 6196 5138 6208
rect 5445 6205 5457 6208
rect 5491 6205 5503 6239
rect 5445 6199 5503 6205
rect 6080 6239 6138 6245
rect 6080 6205 6092 6239
rect 6126 6236 6138 6239
rect 6822 6236 6828 6248
rect 6126 6208 6828 6236
rect 6126 6205 6138 6208
rect 6080 6199 6138 6205
rect 6822 6196 6828 6208
rect 6880 6196 6886 6248
rect 8846 6196 8852 6248
rect 8904 6196 8910 6248
rect 9122 6196 9128 6248
rect 9180 6196 9186 6248
rect 9309 6239 9367 6245
rect 9309 6205 9321 6239
rect 9355 6205 9367 6239
rect 9309 6199 9367 6205
rect 3697 6171 3755 6177
rect 3697 6137 3709 6171
rect 3743 6168 3755 6171
rect 4154 6168 4160 6180
rect 3743 6140 4160 6168
rect 3743 6137 3755 6140
rect 3697 6131 3755 6137
rect 4154 6128 4160 6140
rect 4212 6128 4218 6180
rect 9324 6168 9352 6199
rect 9674 6196 9680 6248
rect 9732 6236 9738 6248
rect 10873 6239 10931 6245
rect 10873 6236 10885 6239
rect 9732 6208 10885 6236
rect 9732 6196 9738 6208
rect 10873 6205 10885 6208
rect 10919 6205 10931 6239
rect 10873 6199 10931 6205
rect 10318 6168 10324 6180
rect 9324 6140 10324 6168
rect 10318 6128 10324 6140
rect 10376 6128 10382 6180
rect 10628 6171 10686 6177
rect 10628 6137 10640 6171
rect 10674 6168 10686 6171
rect 10778 6168 10784 6180
rect 10674 6140 10784 6168
rect 10674 6137 10686 6140
rect 10628 6131 10686 6137
rect 10778 6128 10784 6140
rect 10836 6128 10842 6180
rect 2958 6060 2964 6112
rect 3016 6100 3022 6112
rect 3881 6103 3939 6109
rect 3881 6100 3893 6103
rect 3016 6072 3893 6100
rect 3016 6060 3022 6072
rect 3881 6069 3893 6072
rect 3927 6069 3939 6103
rect 3881 6063 3939 6069
rect 7926 6060 7932 6112
rect 7984 6100 7990 6112
rect 9490 6100 9496 6112
rect 7984 6072 9496 6100
rect 7984 6060 7990 6072
rect 9490 6060 9496 6072
rect 9548 6060 9554 6112
rect 552 6010 11568 6032
rect 552 5958 3112 6010
rect 3164 5958 3176 6010
rect 3228 5958 3240 6010
rect 3292 5958 3304 6010
rect 3356 5958 3368 6010
rect 3420 5958 5826 6010
rect 5878 5958 5890 6010
rect 5942 5958 5954 6010
rect 6006 5958 6018 6010
rect 6070 5958 6082 6010
rect 6134 5958 8540 6010
rect 8592 5958 8604 6010
rect 8656 5958 8668 6010
rect 8720 5958 8732 6010
rect 8784 5958 8796 6010
rect 8848 5958 11254 6010
rect 11306 5958 11318 6010
rect 11370 5958 11382 6010
rect 11434 5958 11446 6010
rect 11498 5958 11510 6010
rect 11562 5958 11568 6010
rect 552 5936 11568 5958
rect 7650 5856 7656 5908
rect 7708 5856 7714 5908
rect 8757 5899 8815 5905
rect 8757 5865 8769 5899
rect 8803 5896 8815 5899
rect 9122 5896 9128 5908
rect 8803 5868 9128 5896
rect 8803 5865 8815 5868
rect 8757 5859 8815 5865
rect 9122 5856 9128 5868
rect 9180 5856 9186 5908
rect 9214 5856 9220 5908
rect 9272 5856 9278 5908
rect 10689 5899 10747 5905
rect 10689 5865 10701 5899
rect 10735 5896 10747 5899
rect 10870 5896 10876 5908
rect 10735 5868 10876 5896
rect 10735 5865 10747 5868
rect 10689 5859 10747 5865
rect 10870 5856 10876 5868
rect 10928 5856 10934 5908
rect 7558 5828 7564 5840
rect 7392 5800 7564 5828
rect 7392 5769 7420 5800
rect 7558 5788 7564 5800
rect 7616 5788 7622 5840
rect 8294 5788 8300 5840
rect 8352 5828 8358 5840
rect 10226 5828 10232 5840
rect 8352 5800 10232 5828
rect 8352 5788 8358 5800
rect 7377 5763 7435 5769
rect 7377 5729 7389 5763
rect 7423 5729 7435 5763
rect 7377 5723 7435 5729
rect 7469 5763 7527 5769
rect 7469 5729 7481 5763
rect 7515 5760 7527 5763
rect 7742 5760 7748 5772
rect 7515 5732 7748 5760
rect 7515 5729 7527 5732
rect 7469 5723 7527 5729
rect 7742 5720 7748 5732
rect 7800 5720 7806 5772
rect 8386 5720 8392 5772
rect 8444 5760 8450 5772
rect 8864 5769 8892 5800
rect 10226 5788 10232 5800
rect 10284 5788 10290 5840
rect 8665 5763 8723 5769
rect 8665 5760 8677 5763
rect 8444 5732 8677 5760
rect 8444 5720 8450 5732
rect 8665 5729 8677 5732
rect 8711 5729 8723 5763
rect 8665 5723 8723 5729
rect 8849 5763 8907 5769
rect 8849 5729 8861 5763
rect 8895 5729 8907 5763
rect 8849 5723 8907 5729
rect 8938 5720 8944 5772
rect 8996 5760 9002 5772
rect 9125 5763 9183 5769
rect 9125 5760 9137 5763
rect 8996 5732 9137 5760
rect 8996 5720 9002 5732
rect 9125 5729 9137 5732
rect 9171 5729 9183 5763
rect 9125 5723 9183 5729
rect 9401 5763 9459 5769
rect 9401 5729 9413 5763
rect 9447 5760 9459 5763
rect 9490 5760 9496 5772
rect 9447 5732 9496 5760
rect 9447 5729 9459 5732
rect 9401 5723 9459 5729
rect 9140 5692 9168 5723
rect 9490 5720 9496 5732
rect 9548 5720 9554 5772
rect 9858 5720 9864 5772
rect 9916 5720 9922 5772
rect 10413 5763 10471 5769
rect 10413 5729 10425 5763
rect 10459 5760 10471 5763
rect 10505 5763 10563 5769
rect 10505 5760 10517 5763
rect 10459 5732 10517 5760
rect 10459 5729 10471 5732
rect 10413 5723 10471 5729
rect 10505 5729 10517 5732
rect 10551 5729 10563 5763
rect 10505 5723 10563 5729
rect 10781 5763 10839 5769
rect 10781 5729 10793 5763
rect 10827 5729 10839 5763
rect 10781 5723 10839 5729
rect 10594 5692 10600 5704
rect 9140 5664 10600 5692
rect 10594 5652 10600 5664
rect 10652 5692 10658 5704
rect 10796 5692 10824 5723
rect 10652 5664 10824 5692
rect 10652 5652 10658 5664
rect 9398 5584 9404 5636
rect 9456 5584 9462 5636
rect 10502 5584 10508 5636
rect 10560 5584 10566 5636
rect 552 5466 11408 5488
rect 552 5414 1755 5466
rect 1807 5414 1819 5466
rect 1871 5414 1883 5466
rect 1935 5414 1947 5466
rect 1999 5414 2011 5466
rect 2063 5414 4469 5466
rect 4521 5414 4533 5466
rect 4585 5414 4597 5466
rect 4649 5414 4661 5466
rect 4713 5414 4725 5466
rect 4777 5414 7183 5466
rect 7235 5414 7247 5466
rect 7299 5414 7311 5466
rect 7363 5414 7375 5466
rect 7427 5414 7439 5466
rect 7491 5414 9897 5466
rect 9949 5414 9961 5466
rect 10013 5414 10025 5466
rect 10077 5414 10089 5466
rect 10141 5414 10153 5466
rect 10205 5414 11408 5466
rect 552 5392 11408 5414
rect 10318 5312 10324 5364
rect 10376 5312 10382 5364
rect 10594 5312 10600 5364
rect 10652 5312 10658 5364
rect 10226 5244 10232 5296
rect 10284 5284 10290 5296
rect 10413 5287 10471 5293
rect 10413 5284 10425 5287
rect 10284 5256 10425 5284
rect 10284 5244 10290 5256
rect 10413 5253 10425 5256
rect 10459 5253 10471 5287
rect 10413 5247 10471 5253
rect 9953 5219 10011 5225
rect 9953 5185 9965 5219
rect 9999 5216 10011 5219
rect 10612 5216 10640 5312
rect 9999 5188 10640 5216
rect 9999 5185 10011 5188
rect 9953 5179 10011 5185
rect 10137 5151 10195 5157
rect 10137 5117 10149 5151
rect 10183 5148 10195 5151
rect 10410 5148 10416 5160
rect 10183 5120 10416 5148
rect 10183 5117 10195 5120
rect 10137 5111 10195 5117
rect 10410 5108 10416 5120
rect 10468 5108 10474 5160
rect 10428 5080 10456 5108
rect 10565 5083 10623 5089
rect 10565 5080 10577 5083
rect 10428 5052 10577 5080
rect 10565 5049 10577 5052
rect 10611 5049 10623 5083
rect 10565 5043 10623 5049
rect 10781 5083 10839 5089
rect 10781 5049 10793 5083
rect 10827 5080 10839 5083
rect 10962 5080 10968 5092
rect 10827 5052 10968 5080
rect 10827 5049 10839 5052
rect 10781 5043 10839 5049
rect 10962 5040 10968 5052
rect 11020 5040 11026 5092
rect 552 4922 11568 4944
rect 552 4870 3112 4922
rect 3164 4870 3176 4922
rect 3228 4870 3240 4922
rect 3292 4870 3304 4922
rect 3356 4870 3368 4922
rect 3420 4870 5826 4922
rect 5878 4870 5890 4922
rect 5942 4870 5954 4922
rect 6006 4870 6018 4922
rect 6070 4870 6082 4922
rect 6134 4870 8540 4922
rect 8592 4870 8604 4922
rect 8656 4870 8668 4922
rect 8720 4870 8732 4922
rect 8784 4870 8796 4922
rect 8848 4870 11254 4922
rect 11306 4870 11318 4922
rect 11370 4870 11382 4922
rect 11434 4870 11446 4922
rect 11498 4870 11510 4922
rect 11562 4870 11568 4922
rect 552 4848 11568 4870
rect 10778 4768 10784 4820
rect 10836 4768 10842 4820
rect 10318 4700 10324 4752
rect 10376 4740 10382 4752
rect 10376 4712 10824 4740
rect 10376 4700 10382 4712
rect 9490 4632 9496 4684
rect 9548 4672 9554 4684
rect 10505 4675 10563 4681
rect 10505 4672 10517 4675
rect 9548 4644 10517 4672
rect 9548 4632 9554 4644
rect 10505 4641 10517 4644
rect 10551 4641 10563 4675
rect 10505 4635 10563 4641
rect 10686 4632 10692 4684
rect 10744 4632 10750 4684
rect 10796 4681 10824 4712
rect 10781 4675 10839 4681
rect 10781 4641 10793 4675
rect 10827 4641 10839 4675
rect 10781 4635 10839 4641
rect 552 4378 11408 4400
rect 552 4326 1755 4378
rect 1807 4326 1819 4378
rect 1871 4326 1883 4378
rect 1935 4326 1947 4378
rect 1999 4326 2011 4378
rect 2063 4326 4469 4378
rect 4521 4326 4533 4378
rect 4585 4326 4597 4378
rect 4649 4326 4661 4378
rect 4713 4326 4725 4378
rect 4777 4326 7183 4378
rect 7235 4326 7247 4378
rect 7299 4326 7311 4378
rect 7363 4326 7375 4378
rect 7427 4326 7439 4378
rect 7491 4326 9897 4378
rect 9949 4326 9961 4378
rect 10013 4326 10025 4378
rect 10077 4326 10089 4378
rect 10141 4326 10153 4378
rect 10205 4326 11408 4378
rect 552 4304 11408 4326
rect 552 3834 11568 3856
rect 552 3782 3112 3834
rect 3164 3782 3176 3834
rect 3228 3782 3240 3834
rect 3292 3782 3304 3834
rect 3356 3782 3368 3834
rect 3420 3782 5826 3834
rect 5878 3782 5890 3834
rect 5942 3782 5954 3834
rect 6006 3782 6018 3834
rect 6070 3782 6082 3834
rect 6134 3782 8540 3834
rect 8592 3782 8604 3834
rect 8656 3782 8668 3834
rect 8720 3782 8732 3834
rect 8784 3782 8796 3834
rect 8848 3782 11254 3834
rect 11306 3782 11318 3834
rect 11370 3782 11382 3834
rect 11434 3782 11446 3834
rect 11498 3782 11510 3834
rect 11562 3782 11568 3834
rect 552 3760 11568 3782
rect 552 3290 11408 3312
rect 552 3238 1755 3290
rect 1807 3238 1819 3290
rect 1871 3238 1883 3290
rect 1935 3238 1947 3290
rect 1999 3238 2011 3290
rect 2063 3238 4469 3290
rect 4521 3238 4533 3290
rect 4585 3238 4597 3290
rect 4649 3238 4661 3290
rect 4713 3238 4725 3290
rect 4777 3238 7183 3290
rect 7235 3238 7247 3290
rect 7299 3238 7311 3290
rect 7363 3238 7375 3290
rect 7427 3238 7439 3290
rect 7491 3238 9897 3290
rect 9949 3238 9961 3290
rect 10013 3238 10025 3290
rect 10077 3238 10089 3290
rect 10141 3238 10153 3290
rect 10205 3238 11408 3290
rect 552 3216 11408 3238
rect 552 2746 11568 2768
rect 552 2694 3112 2746
rect 3164 2694 3176 2746
rect 3228 2694 3240 2746
rect 3292 2694 3304 2746
rect 3356 2694 3368 2746
rect 3420 2694 5826 2746
rect 5878 2694 5890 2746
rect 5942 2694 5954 2746
rect 6006 2694 6018 2746
rect 6070 2694 6082 2746
rect 6134 2694 8540 2746
rect 8592 2694 8604 2746
rect 8656 2694 8668 2746
rect 8720 2694 8732 2746
rect 8784 2694 8796 2746
rect 8848 2694 11254 2746
rect 11306 2694 11318 2746
rect 11370 2694 11382 2746
rect 11434 2694 11446 2746
rect 11498 2694 11510 2746
rect 11562 2694 11568 2746
rect 552 2672 11568 2694
rect 552 2202 11408 2224
rect 552 2150 1755 2202
rect 1807 2150 1819 2202
rect 1871 2150 1883 2202
rect 1935 2150 1947 2202
rect 1999 2150 2011 2202
rect 2063 2150 4469 2202
rect 4521 2150 4533 2202
rect 4585 2150 4597 2202
rect 4649 2150 4661 2202
rect 4713 2150 4725 2202
rect 4777 2150 7183 2202
rect 7235 2150 7247 2202
rect 7299 2150 7311 2202
rect 7363 2150 7375 2202
rect 7427 2150 7439 2202
rect 7491 2150 9897 2202
rect 9949 2150 9961 2202
rect 10013 2150 10025 2202
rect 10077 2150 10089 2202
rect 10141 2150 10153 2202
rect 10205 2150 11408 2202
rect 552 2128 11408 2150
rect 552 1658 11568 1680
rect 552 1606 3112 1658
rect 3164 1606 3176 1658
rect 3228 1606 3240 1658
rect 3292 1606 3304 1658
rect 3356 1606 3368 1658
rect 3420 1606 5826 1658
rect 5878 1606 5890 1658
rect 5942 1606 5954 1658
rect 6006 1606 6018 1658
rect 6070 1606 6082 1658
rect 6134 1606 8540 1658
rect 8592 1606 8604 1658
rect 8656 1606 8668 1658
rect 8720 1606 8732 1658
rect 8784 1606 8796 1658
rect 8848 1606 11254 1658
rect 11306 1606 11318 1658
rect 11370 1606 11382 1658
rect 11434 1606 11446 1658
rect 11498 1606 11510 1658
rect 11562 1606 11568 1658
rect 552 1584 11568 1606
rect 552 1114 11408 1136
rect 552 1062 1755 1114
rect 1807 1062 1819 1114
rect 1871 1062 1883 1114
rect 1935 1062 1947 1114
rect 1999 1062 2011 1114
rect 2063 1062 4469 1114
rect 4521 1062 4533 1114
rect 4585 1062 4597 1114
rect 4649 1062 4661 1114
rect 4713 1062 4725 1114
rect 4777 1062 7183 1114
rect 7235 1062 7247 1114
rect 7299 1062 7311 1114
rect 7363 1062 7375 1114
rect 7427 1062 7439 1114
rect 7491 1062 9897 1114
rect 9949 1062 9961 1114
rect 10013 1062 10025 1114
rect 10077 1062 10089 1114
rect 10141 1062 10153 1114
rect 10205 1062 11408 1114
rect 552 1040 11408 1062
rect 552 570 11568 592
rect 552 518 3112 570
rect 3164 518 3176 570
rect 3228 518 3240 570
rect 3292 518 3304 570
rect 3356 518 3368 570
rect 3420 518 5826 570
rect 5878 518 5890 570
rect 5942 518 5954 570
rect 6006 518 6018 570
rect 6070 518 6082 570
rect 6134 518 8540 570
rect 8592 518 8604 570
rect 8656 518 8668 570
rect 8720 518 8732 570
rect 8784 518 8796 570
rect 8848 518 11254 570
rect 11306 518 11318 570
rect 11370 518 11382 570
rect 11434 518 11446 570
rect 11498 518 11510 570
rect 11562 518 11568 570
rect 552 496 11568 518
<< via1 >>
rect 3976 11636 4028 11688
rect 7840 11636 7892 11688
rect 9588 11636 9640 11688
rect 6644 11568 6696 11620
rect 8024 11568 8076 11620
rect 8300 11568 8352 11620
rect 8484 11568 8536 11620
rect 2872 11500 2924 11552
rect 3332 11500 3384 11552
rect 5908 11500 5960 11552
rect 6184 11500 6236 11552
rect 7196 11500 7248 11552
rect 9496 11500 9548 11552
rect 3112 11398 3164 11450
rect 3176 11398 3228 11450
rect 3240 11398 3292 11450
rect 3304 11398 3356 11450
rect 3368 11398 3420 11450
rect 5826 11398 5878 11450
rect 5890 11398 5942 11450
rect 5954 11398 6006 11450
rect 6018 11398 6070 11450
rect 6082 11398 6134 11450
rect 8540 11398 8592 11450
rect 8604 11398 8656 11450
rect 8668 11398 8720 11450
rect 8732 11398 8784 11450
rect 8796 11398 8848 11450
rect 11254 11398 11306 11450
rect 11318 11398 11370 11450
rect 11382 11398 11434 11450
rect 11446 11398 11498 11450
rect 11510 11398 11562 11450
rect 4620 11296 4672 11348
rect 6184 11296 6236 11348
rect 8300 11296 8352 11348
rect 2688 11271 2740 11280
rect 2688 11237 2697 11271
rect 2697 11237 2731 11271
rect 2731 11237 2740 11271
rect 2688 11228 2740 11237
rect 3976 11228 4028 11280
rect 3056 11160 3108 11212
rect 5172 11203 5224 11212
rect 5172 11169 5181 11203
rect 5181 11169 5215 11203
rect 5215 11169 5224 11203
rect 5172 11160 5224 11169
rect 3608 11135 3660 11144
rect 3608 11101 3617 11135
rect 3617 11101 3651 11135
rect 3651 11101 3660 11135
rect 3608 11092 3660 11101
rect 3792 11092 3844 11144
rect 6644 11203 6696 11212
rect 6644 11169 6653 11203
rect 6653 11169 6687 11203
rect 6687 11169 6696 11203
rect 6644 11160 6696 11169
rect 7656 11228 7708 11280
rect 7104 11160 7156 11212
rect 7564 11203 7616 11212
rect 7564 11169 7573 11203
rect 7573 11169 7607 11203
rect 7607 11169 7616 11203
rect 7564 11160 7616 11169
rect 7840 11160 7892 11212
rect 8024 11203 8076 11212
rect 8024 11169 8033 11203
rect 8033 11169 8067 11203
rect 8067 11169 8076 11203
rect 8024 11160 8076 11169
rect 11060 11228 11112 11280
rect 8944 11160 8996 11212
rect 6920 11092 6972 11144
rect 7012 11092 7064 11144
rect 7196 11135 7248 11144
rect 7196 11101 7205 11135
rect 7205 11101 7239 11135
rect 7239 11101 7248 11135
rect 7196 11092 7248 11101
rect 8116 11092 8168 11144
rect 5540 11024 5592 11076
rect 7288 11024 7340 11076
rect 7656 11024 7708 11076
rect 7932 11024 7984 11076
rect 2964 10956 3016 11008
rect 3700 10956 3752 11008
rect 4988 10999 5040 11008
rect 4988 10965 4997 10999
rect 4997 10965 5031 10999
rect 5031 10965 5040 10999
rect 4988 10956 5040 10965
rect 6736 10956 6788 11008
rect 7564 10999 7616 11008
rect 7564 10965 7573 10999
rect 7573 10965 7607 10999
rect 7607 10965 7616 10999
rect 7564 10956 7616 10965
rect 7748 10956 7800 11008
rect 10784 11135 10836 11144
rect 10784 11101 10793 11135
rect 10793 11101 10827 11135
rect 10827 11101 10836 11135
rect 10784 11092 10836 11101
rect 10232 10956 10284 11008
rect 1755 10854 1807 10906
rect 1819 10854 1871 10906
rect 1883 10854 1935 10906
rect 1947 10854 1999 10906
rect 2011 10854 2063 10906
rect 4469 10854 4521 10906
rect 4533 10854 4585 10906
rect 4597 10854 4649 10906
rect 4661 10854 4713 10906
rect 4725 10854 4777 10906
rect 7183 10854 7235 10906
rect 7247 10854 7299 10906
rect 7311 10854 7363 10906
rect 7375 10854 7427 10906
rect 7439 10854 7491 10906
rect 9897 10854 9949 10906
rect 9961 10854 10013 10906
rect 10025 10854 10077 10906
rect 10089 10854 10141 10906
rect 10153 10854 10205 10906
rect 756 10752 808 10804
rect 2136 10752 2188 10804
rect 2872 10795 2924 10804
rect 2872 10761 2881 10795
rect 2881 10761 2915 10795
rect 2915 10761 2924 10795
rect 2872 10752 2924 10761
rect 3056 10752 3108 10804
rect 6736 10752 6788 10804
rect 1032 10684 1084 10736
rect 3792 10684 3844 10736
rect 4068 10684 4120 10736
rect 6920 10684 6972 10736
rect 1308 10548 1360 10600
rect 1676 10548 1728 10600
rect 3056 10591 3108 10600
rect 3056 10557 3065 10591
rect 3065 10557 3099 10591
rect 3099 10557 3108 10591
rect 3056 10548 3108 10557
rect 3240 10591 3292 10600
rect 3240 10557 3249 10591
rect 3249 10557 3283 10591
rect 3283 10557 3292 10591
rect 3240 10548 3292 10557
rect 3608 10548 3660 10600
rect 3700 10548 3752 10600
rect 3976 10591 4028 10600
rect 3976 10557 3985 10591
rect 3985 10557 4019 10591
rect 4019 10557 4028 10591
rect 3976 10548 4028 10557
rect 4160 10548 4212 10600
rect 8300 10752 8352 10804
rect 8208 10727 8260 10736
rect 8208 10693 8217 10727
rect 8217 10693 8251 10727
rect 8251 10693 8260 10727
rect 8208 10684 8260 10693
rect 1216 10480 1268 10532
rect 2596 10455 2648 10464
rect 2596 10421 2605 10455
rect 2605 10421 2639 10455
rect 2639 10421 2648 10455
rect 2596 10412 2648 10421
rect 4804 10480 4856 10532
rect 7472 10548 7524 10600
rect 7748 10548 7800 10600
rect 8024 10616 8076 10668
rect 10784 10659 10836 10668
rect 10784 10625 10793 10659
rect 10793 10625 10827 10659
rect 10827 10625 10836 10659
rect 10784 10616 10836 10625
rect 5356 10480 5408 10532
rect 5724 10480 5776 10532
rect 11060 10591 11112 10600
rect 11060 10557 11069 10591
rect 11069 10557 11103 10591
rect 11103 10557 11112 10591
rect 11060 10548 11112 10557
rect 6736 10455 6788 10464
rect 6736 10421 6745 10455
rect 6745 10421 6779 10455
rect 6779 10421 6788 10455
rect 6736 10412 6788 10421
rect 7104 10412 7156 10464
rect 7932 10412 7984 10464
rect 9312 10455 9364 10464
rect 9312 10421 9321 10455
rect 9321 10421 9355 10455
rect 9355 10421 9364 10455
rect 9312 10412 9364 10421
rect 3112 10310 3164 10362
rect 3176 10310 3228 10362
rect 3240 10310 3292 10362
rect 3304 10310 3356 10362
rect 3368 10310 3420 10362
rect 5826 10310 5878 10362
rect 5890 10310 5942 10362
rect 5954 10310 6006 10362
rect 6018 10310 6070 10362
rect 6082 10310 6134 10362
rect 8540 10310 8592 10362
rect 8604 10310 8656 10362
rect 8668 10310 8720 10362
rect 8732 10310 8784 10362
rect 8796 10310 8848 10362
rect 11254 10310 11306 10362
rect 11318 10310 11370 10362
rect 11382 10310 11434 10362
rect 11446 10310 11498 10362
rect 11510 10310 11562 10362
rect 1124 10140 1176 10192
rect 1032 10115 1084 10124
rect 1032 10081 1041 10115
rect 1041 10081 1075 10115
rect 1075 10081 1084 10115
rect 1032 10072 1084 10081
rect 1216 10115 1268 10124
rect 1216 10081 1225 10115
rect 1225 10081 1259 10115
rect 1259 10081 1268 10115
rect 1216 10072 1268 10081
rect 2688 10208 2740 10260
rect 2872 10140 2924 10192
rect 2412 10072 2464 10124
rect 2780 10115 2832 10124
rect 3516 10208 3568 10260
rect 3700 10208 3752 10260
rect 4988 10140 5040 10192
rect 2780 10081 2798 10115
rect 2798 10081 2832 10115
rect 2780 10072 2832 10081
rect 3424 10072 3476 10124
rect 4160 10072 4212 10124
rect 5356 10208 5408 10260
rect 3056 10047 3108 10056
rect 3056 10013 3065 10047
rect 3065 10013 3099 10047
rect 3099 10013 3108 10047
rect 3056 10004 3108 10013
rect 4804 10047 4856 10056
rect 4804 10013 4813 10047
rect 4813 10013 4847 10047
rect 4847 10013 4856 10047
rect 4804 10004 4856 10013
rect 5540 10115 5592 10124
rect 5540 10081 5549 10115
rect 5549 10081 5583 10115
rect 5583 10081 5592 10115
rect 5540 10072 5592 10081
rect 6736 10140 6788 10192
rect 7564 10208 7616 10260
rect 8116 10208 8168 10260
rect 9496 10251 9548 10260
rect 9496 10217 9505 10251
rect 9505 10217 9539 10251
rect 9539 10217 9548 10251
rect 9496 10208 9548 10217
rect 9588 10208 9640 10260
rect 7012 10115 7064 10124
rect 7012 10081 7021 10115
rect 7021 10081 7055 10115
rect 7055 10081 7064 10115
rect 7012 10072 7064 10081
rect 9680 10140 9732 10192
rect 7656 10072 7708 10124
rect 7840 10072 7892 10124
rect 8208 10072 8260 10124
rect 1676 9979 1728 9988
rect 1676 9945 1685 9979
rect 1685 9945 1719 9979
rect 1719 9945 1728 9979
rect 1676 9936 1728 9945
rect 7104 9936 7156 9988
rect 8300 9936 8352 9988
rect 10508 10047 10560 10056
rect 10508 10013 10517 10047
rect 10517 10013 10551 10047
rect 10551 10013 10560 10047
rect 10508 10004 10560 10013
rect 1216 9911 1268 9920
rect 1216 9877 1225 9911
rect 1225 9877 1259 9911
rect 1259 9877 1268 9911
rect 1216 9868 1268 9877
rect 1584 9911 1636 9920
rect 1584 9877 1593 9911
rect 1593 9877 1627 9911
rect 1627 9877 1636 9911
rect 1584 9868 1636 9877
rect 3608 9868 3660 9920
rect 3884 9868 3936 9920
rect 5816 9911 5868 9920
rect 5816 9877 5825 9911
rect 5825 9877 5859 9911
rect 5859 9877 5868 9911
rect 5816 9868 5868 9877
rect 7012 9868 7064 9920
rect 7748 9868 7800 9920
rect 8024 9868 8076 9920
rect 9772 9868 9824 9920
rect 1755 9766 1807 9818
rect 1819 9766 1871 9818
rect 1883 9766 1935 9818
rect 1947 9766 1999 9818
rect 2011 9766 2063 9818
rect 4469 9766 4521 9818
rect 4533 9766 4585 9818
rect 4597 9766 4649 9818
rect 4661 9766 4713 9818
rect 4725 9766 4777 9818
rect 7183 9766 7235 9818
rect 7247 9766 7299 9818
rect 7311 9766 7363 9818
rect 7375 9766 7427 9818
rect 7439 9766 7491 9818
rect 9897 9766 9949 9818
rect 9961 9766 10013 9818
rect 10025 9766 10077 9818
rect 10089 9766 10141 9818
rect 10153 9766 10205 9818
rect 1308 9707 1360 9716
rect 1308 9673 1317 9707
rect 1317 9673 1351 9707
rect 1351 9673 1360 9707
rect 1308 9664 1360 9673
rect 1124 9639 1176 9648
rect 1124 9605 1133 9639
rect 1133 9605 1167 9639
rect 1167 9605 1176 9639
rect 1124 9596 1176 9605
rect 3056 9596 3108 9648
rect 4896 9596 4948 9648
rect 5448 9596 5500 9648
rect 7012 9707 7064 9716
rect 7012 9673 7021 9707
rect 7021 9673 7055 9707
rect 7055 9673 7064 9707
rect 7012 9664 7064 9673
rect 8208 9664 8260 9716
rect 8944 9664 8996 9716
rect 7288 9596 7340 9648
rect 1584 9460 1636 9512
rect 3056 9503 3108 9512
rect 3056 9469 3065 9503
rect 3065 9469 3099 9503
rect 3099 9469 3108 9503
rect 3056 9460 3108 9469
rect 3516 9460 3568 9512
rect 4804 9528 4856 9580
rect 7748 9528 7800 9580
rect 5448 9460 5500 9512
rect 8300 9596 8352 9648
rect 10600 9596 10652 9648
rect 3332 9392 3384 9444
rect 4896 9392 4948 9444
rect 5264 9435 5316 9444
rect 5264 9401 5273 9435
rect 5273 9401 5307 9435
rect 5307 9401 5316 9435
rect 5264 9392 5316 9401
rect 5908 9435 5960 9444
rect 5908 9401 5942 9435
rect 5942 9401 5960 9435
rect 5908 9392 5960 9401
rect 2596 9324 2648 9376
rect 4068 9324 4120 9376
rect 7104 9367 7156 9376
rect 7104 9333 7113 9367
rect 7113 9333 7147 9367
rect 7147 9333 7156 9367
rect 7104 9324 7156 9333
rect 7288 9367 7340 9376
rect 7288 9333 7297 9367
rect 7297 9333 7331 9367
rect 7331 9333 7340 9367
rect 7288 9324 7340 9333
rect 7564 9392 7616 9444
rect 8116 9435 8168 9444
rect 8116 9401 8125 9435
rect 8125 9401 8159 9435
rect 8159 9401 8168 9435
rect 8116 9392 8168 9401
rect 7748 9367 7800 9376
rect 7748 9333 7757 9367
rect 7757 9333 7791 9367
rect 7791 9333 7800 9367
rect 7748 9324 7800 9333
rect 8024 9324 8076 9376
rect 8668 9503 8720 9512
rect 8668 9469 8677 9503
rect 8677 9469 8711 9503
rect 8711 9469 8720 9503
rect 8668 9460 8720 9469
rect 9680 9460 9732 9512
rect 10324 9460 10376 9512
rect 9036 9392 9088 9444
rect 10232 9324 10284 9376
rect 10416 9367 10468 9376
rect 10416 9333 10425 9367
rect 10425 9333 10459 9367
rect 10459 9333 10468 9367
rect 10416 9324 10468 9333
rect 3112 9222 3164 9274
rect 3176 9222 3228 9274
rect 3240 9222 3292 9274
rect 3304 9222 3356 9274
rect 3368 9222 3420 9274
rect 5826 9222 5878 9274
rect 5890 9222 5942 9274
rect 5954 9222 6006 9274
rect 6018 9222 6070 9274
rect 6082 9222 6134 9274
rect 8540 9222 8592 9274
rect 8604 9222 8656 9274
rect 8668 9222 8720 9274
rect 8732 9222 8784 9274
rect 8796 9222 8848 9274
rect 11254 9222 11306 9274
rect 11318 9222 11370 9274
rect 11382 9222 11434 9274
rect 11446 9222 11498 9274
rect 11510 9222 11562 9274
rect 2412 9163 2464 9172
rect 2412 9129 2421 9163
rect 2421 9129 2455 9163
rect 2455 9129 2464 9163
rect 2412 9120 2464 9129
rect 2872 9120 2924 9172
rect 3792 9120 3844 9172
rect 5724 9120 5776 9172
rect 3976 9052 4028 9104
rect 9036 9120 9088 9172
rect 10324 9095 10376 9104
rect 10324 9061 10333 9095
rect 10333 9061 10367 9095
rect 10367 9061 10376 9095
rect 10324 9052 10376 9061
rect 11060 9052 11112 9104
rect 4160 8984 4212 9036
rect 6368 8984 6420 9036
rect 7840 9027 7892 9036
rect 7840 8993 7849 9027
rect 7849 8993 7883 9027
rect 7883 8993 7892 9027
rect 7840 8984 7892 8993
rect 2596 8848 2648 8900
rect 3700 8959 3752 8968
rect 3700 8925 3709 8959
rect 3709 8925 3743 8959
rect 3743 8925 3752 8959
rect 3700 8916 3752 8925
rect 5448 8916 5500 8968
rect 7932 8916 7984 8968
rect 10416 8984 10468 9036
rect 9772 8916 9824 8968
rect 10232 8916 10284 8968
rect 10784 8959 10836 8968
rect 10784 8925 10793 8959
rect 10793 8925 10827 8959
rect 10827 8925 10836 8959
rect 10784 8916 10836 8925
rect 3332 8780 3384 8832
rect 4068 8780 4120 8832
rect 7656 8780 7708 8832
rect 8116 8780 8168 8832
rect 8300 8780 8352 8832
rect 10416 8823 10468 8832
rect 10416 8789 10425 8823
rect 10425 8789 10459 8823
rect 10459 8789 10468 8823
rect 10416 8780 10468 8789
rect 1755 8678 1807 8730
rect 1819 8678 1871 8730
rect 1883 8678 1935 8730
rect 1947 8678 1999 8730
rect 2011 8678 2063 8730
rect 4469 8678 4521 8730
rect 4533 8678 4585 8730
rect 4597 8678 4649 8730
rect 4661 8678 4713 8730
rect 4725 8678 4777 8730
rect 7183 8678 7235 8730
rect 7247 8678 7299 8730
rect 7311 8678 7363 8730
rect 7375 8678 7427 8730
rect 7439 8678 7491 8730
rect 9897 8678 9949 8730
rect 9961 8678 10013 8730
rect 10025 8678 10077 8730
rect 10089 8678 10141 8730
rect 10153 8678 10205 8730
rect 2780 8576 2832 8628
rect 2964 8372 3016 8424
rect 7012 8576 7064 8628
rect 3516 8508 3568 8560
rect 4068 8508 4120 8560
rect 5172 8508 5224 8560
rect 2964 8236 3016 8288
rect 3608 8372 3660 8424
rect 4712 8440 4764 8492
rect 3332 8304 3384 8356
rect 3976 8415 4028 8424
rect 3976 8381 3985 8415
rect 3985 8381 4019 8415
rect 4019 8381 4028 8415
rect 3976 8372 4028 8381
rect 7748 8576 7800 8628
rect 4160 8347 4212 8356
rect 4160 8313 4169 8347
rect 4169 8313 4203 8347
rect 4203 8313 4212 8347
rect 4160 8304 4212 8313
rect 4804 8304 4856 8356
rect 5724 8372 5776 8424
rect 7104 8440 7156 8492
rect 6276 8372 6328 8424
rect 6460 8415 6512 8424
rect 6460 8381 6469 8415
rect 6469 8381 6503 8415
rect 6503 8381 6512 8415
rect 6460 8372 6512 8381
rect 4988 8347 5040 8356
rect 4988 8313 4997 8347
rect 4997 8313 5031 8347
rect 5031 8313 5040 8347
rect 4988 8304 5040 8313
rect 5080 8304 5132 8356
rect 6644 8304 6696 8356
rect 6828 8415 6880 8424
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 6920 8415 6972 8424
rect 6920 8381 6929 8415
rect 6929 8381 6963 8415
rect 6963 8381 6972 8415
rect 6920 8372 6972 8381
rect 7196 8415 7248 8424
rect 7196 8381 7205 8415
rect 7205 8381 7239 8415
rect 7239 8381 7248 8415
rect 7196 8372 7248 8381
rect 7472 8372 7524 8424
rect 7748 8372 7800 8424
rect 7932 8415 7984 8424
rect 7932 8381 7941 8415
rect 7941 8381 7975 8415
rect 7975 8381 7984 8415
rect 7932 8372 7984 8381
rect 8208 8415 8260 8424
rect 8208 8381 8217 8415
rect 8217 8381 8251 8415
rect 8251 8381 8260 8415
rect 8208 8372 8260 8381
rect 8392 8347 8444 8356
rect 8392 8313 8401 8347
rect 8401 8313 8435 8347
rect 8435 8313 8444 8347
rect 8392 8304 8444 8313
rect 3792 8279 3844 8288
rect 3792 8245 3801 8279
rect 3801 8245 3835 8279
rect 3835 8245 3844 8279
rect 3792 8236 3844 8245
rect 5172 8279 5224 8288
rect 5172 8245 5181 8279
rect 5181 8245 5215 8279
rect 5215 8245 5224 8279
rect 5172 8236 5224 8245
rect 5264 8279 5316 8288
rect 5264 8245 5273 8279
rect 5273 8245 5307 8279
rect 5307 8245 5316 8279
rect 5264 8236 5316 8245
rect 6184 8236 6236 8288
rect 6828 8236 6880 8288
rect 8852 8415 8904 8424
rect 8852 8381 8861 8415
rect 8861 8381 8895 8415
rect 8895 8381 8904 8415
rect 8852 8372 8904 8381
rect 9680 8372 9732 8424
rect 10324 8372 10376 8424
rect 10968 8415 11020 8424
rect 10968 8381 10977 8415
rect 10977 8381 11011 8415
rect 11011 8381 11020 8415
rect 10968 8372 11020 8381
rect 9036 8304 9088 8356
rect 9496 8304 9548 8356
rect 9312 8236 9364 8288
rect 10968 8236 11020 8288
rect 3112 8134 3164 8186
rect 3176 8134 3228 8186
rect 3240 8134 3292 8186
rect 3304 8134 3356 8186
rect 3368 8134 3420 8186
rect 5826 8134 5878 8186
rect 5890 8134 5942 8186
rect 5954 8134 6006 8186
rect 6018 8134 6070 8186
rect 6082 8134 6134 8186
rect 8540 8134 8592 8186
rect 8604 8134 8656 8186
rect 8668 8134 8720 8186
rect 8732 8134 8784 8186
rect 8796 8134 8848 8186
rect 11254 8134 11306 8186
rect 11318 8134 11370 8186
rect 11382 8134 11434 8186
rect 11446 8134 11498 8186
rect 11510 8134 11562 8186
rect 4712 8032 4764 8084
rect 6460 8032 6512 8084
rect 6920 8032 6972 8084
rect 7564 8032 7616 8084
rect 8116 8032 8168 8084
rect 8944 8075 8996 8084
rect 8944 8041 8953 8075
rect 8953 8041 8987 8075
rect 8987 8041 8996 8075
rect 8944 8032 8996 8041
rect 10508 8032 10560 8084
rect 10600 8075 10652 8084
rect 10600 8041 10609 8075
rect 10609 8041 10643 8075
rect 10643 8041 10652 8075
rect 10600 8032 10652 8041
rect 2780 7939 2832 7948
rect 2780 7905 2789 7939
rect 2789 7905 2823 7939
rect 2823 7905 2832 7939
rect 2780 7896 2832 7905
rect 2964 7896 3016 7948
rect 3700 7964 3752 8016
rect 7656 7964 7708 8016
rect 8024 7964 8076 8016
rect 3424 7939 3476 7948
rect 3424 7905 3458 7939
rect 3458 7905 3476 7939
rect 3424 7896 3476 7905
rect 5264 7896 5316 7948
rect 7564 7896 7616 7948
rect 5448 7871 5500 7880
rect 5448 7837 5457 7871
rect 5457 7837 5491 7871
rect 5491 7837 5500 7871
rect 5448 7828 5500 7837
rect 7196 7828 7248 7880
rect 7472 7828 7524 7880
rect 8208 7828 8260 7880
rect 8944 7896 8996 7948
rect 9404 7896 9456 7948
rect 10416 8007 10468 8016
rect 10416 7973 10425 8007
rect 10425 7973 10459 8007
rect 10459 7973 10468 8007
rect 10416 7964 10468 7973
rect 9128 7828 9180 7880
rect 9772 7828 9824 7880
rect 7748 7760 7800 7812
rect 11152 7828 11204 7880
rect 2596 7735 2648 7744
rect 2596 7701 2605 7735
rect 2605 7701 2639 7735
rect 2639 7701 2648 7735
rect 2596 7692 2648 7701
rect 2964 7735 3016 7744
rect 2964 7701 2973 7735
rect 2973 7701 3007 7735
rect 3007 7701 3016 7735
rect 2964 7692 3016 7701
rect 3332 7692 3384 7744
rect 4988 7692 5040 7744
rect 5356 7692 5408 7744
rect 5540 7692 5592 7744
rect 6368 7692 6420 7744
rect 10968 7760 11020 7812
rect 9220 7692 9272 7744
rect 9588 7692 9640 7744
rect 1755 7590 1807 7642
rect 1819 7590 1871 7642
rect 1883 7590 1935 7642
rect 1947 7590 1999 7642
rect 2011 7590 2063 7642
rect 4469 7590 4521 7642
rect 4533 7590 4585 7642
rect 4597 7590 4649 7642
rect 4661 7590 4713 7642
rect 4725 7590 4777 7642
rect 7183 7590 7235 7642
rect 7247 7590 7299 7642
rect 7311 7590 7363 7642
rect 7375 7590 7427 7642
rect 7439 7590 7491 7642
rect 9897 7590 9949 7642
rect 9961 7590 10013 7642
rect 10025 7590 10077 7642
rect 10089 7590 10141 7642
rect 10153 7590 10205 7642
rect 2964 7488 3016 7540
rect 2596 7352 2648 7404
rect 3516 7488 3568 7540
rect 5172 7488 5224 7540
rect 5448 7531 5500 7540
rect 5448 7497 5457 7531
rect 5457 7497 5491 7531
rect 5491 7497 5500 7531
rect 5448 7488 5500 7497
rect 7104 7488 7156 7540
rect 7932 7488 7984 7540
rect 8208 7531 8260 7540
rect 8208 7497 8217 7531
rect 8217 7497 8251 7531
rect 8251 7497 8260 7531
rect 8208 7488 8260 7497
rect 9312 7531 9364 7540
rect 9312 7497 9321 7531
rect 9321 7497 9355 7531
rect 9355 7497 9364 7531
rect 9312 7488 9364 7497
rect 9220 7395 9272 7404
rect 9220 7361 9229 7395
rect 9229 7361 9263 7395
rect 9263 7361 9272 7395
rect 9220 7352 9272 7361
rect 10784 7352 10836 7404
rect 3700 7327 3752 7336
rect 3700 7293 3709 7327
rect 3709 7293 3743 7327
rect 3743 7293 3752 7327
rect 3700 7284 3752 7293
rect 3792 7284 3844 7336
rect 5172 7327 5224 7336
rect 5172 7293 5181 7327
rect 5181 7293 5215 7327
rect 5215 7293 5224 7327
rect 5172 7284 5224 7293
rect 5264 7284 5316 7336
rect 5540 7284 5592 7336
rect 5632 7327 5684 7336
rect 5632 7293 5641 7327
rect 5641 7293 5675 7327
rect 5675 7293 5684 7327
rect 5632 7284 5684 7293
rect 6184 7284 6236 7336
rect 7104 7327 7156 7336
rect 7104 7293 7113 7327
rect 7113 7293 7147 7327
rect 7147 7293 7156 7327
rect 7104 7284 7156 7293
rect 7748 7284 7800 7336
rect 8944 7327 8996 7336
rect 8944 7293 8953 7327
rect 8953 7293 8987 7327
rect 8987 7293 8996 7327
rect 8944 7284 8996 7293
rect 2504 7216 2556 7268
rect 2964 7216 3016 7268
rect 3332 7216 3384 7268
rect 3608 7191 3660 7200
rect 3608 7157 3617 7191
rect 3617 7157 3651 7191
rect 3651 7157 3660 7191
rect 3608 7148 3660 7157
rect 6736 7216 6788 7268
rect 7932 7216 7984 7268
rect 8208 7216 8260 7268
rect 10508 7284 10560 7336
rect 5356 7148 5408 7200
rect 8116 7148 8168 7200
rect 9220 7148 9272 7200
rect 9772 7148 9824 7200
rect 10692 7148 10744 7200
rect 3112 7046 3164 7098
rect 3176 7046 3228 7098
rect 3240 7046 3292 7098
rect 3304 7046 3356 7098
rect 3368 7046 3420 7098
rect 5826 7046 5878 7098
rect 5890 7046 5942 7098
rect 5954 7046 6006 7098
rect 6018 7046 6070 7098
rect 6082 7046 6134 7098
rect 8540 7046 8592 7098
rect 8604 7046 8656 7098
rect 8668 7046 8720 7098
rect 8732 7046 8784 7098
rect 8796 7046 8848 7098
rect 11254 7046 11306 7098
rect 11318 7046 11370 7098
rect 11382 7046 11434 7098
rect 11446 7046 11498 7098
rect 11510 7046 11562 7098
rect 3516 6944 3568 6996
rect 9128 6944 9180 6996
rect 10784 6944 10836 6996
rect 2504 6851 2556 6860
rect 2504 6817 2538 6851
rect 2538 6817 2556 6851
rect 5632 6876 5684 6928
rect 2504 6808 2556 6817
rect 3700 6783 3752 6792
rect 3700 6749 3709 6783
rect 3709 6749 3743 6783
rect 3743 6749 3752 6783
rect 3976 6851 4028 6860
rect 3976 6817 4010 6851
rect 4010 6817 4028 6851
rect 3976 6808 4028 6817
rect 4252 6808 4304 6860
rect 5724 6808 5776 6860
rect 6092 6851 6144 6860
rect 6092 6817 6101 6851
rect 6101 6817 6135 6851
rect 6135 6817 6144 6851
rect 6092 6808 6144 6817
rect 7104 6876 7156 6928
rect 6644 6851 6696 6860
rect 6644 6817 6678 6851
rect 6678 6817 6696 6851
rect 6644 6808 6696 6817
rect 8392 6808 8444 6860
rect 9588 6851 9640 6860
rect 9588 6817 9622 6851
rect 9622 6817 9640 6851
rect 9588 6808 9640 6817
rect 3700 6740 3752 6749
rect 5080 6715 5132 6724
rect 5080 6681 5089 6715
rect 5089 6681 5123 6715
rect 5123 6681 5132 6715
rect 5080 6672 5132 6681
rect 6276 6715 6328 6724
rect 6276 6681 6285 6715
rect 6285 6681 6319 6715
rect 6319 6681 6328 6715
rect 6276 6672 6328 6681
rect 5356 6647 5408 6656
rect 5356 6613 5365 6647
rect 5365 6613 5399 6647
rect 5399 6613 5408 6647
rect 5356 6604 5408 6613
rect 7748 6647 7800 6656
rect 7748 6613 7757 6647
rect 7757 6613 7791 6647
rect 7791 6613 7800 6647
rect 7748 6604 7800 6613
rect 9680 6604 9732 6656
rect 1755 6502 1807 6554
rect 1819 6502 1871 6554
rect 1883 6502 1935 6554
rect 1947 6502 1999 6554
rect 2011 6502 2063 6554
rect 4469 6502 4521 6554
rect 4533 6502 4585 6554
rect 4597 6502 4649 6554
rect 4661 6502 4713 6554
rect 4725 6502 4777 6554
rect 7183 6502 7235 6554
rect 7247 6502 7299 6554
rect 7311 6502 7363 6554
rect 7375 6502 7427 6554
rect 7439 6502 7491 6554
rect 9897 6502 9949 6554
rect 9961 6502 10013 6554
rect 10025 6502 10077 6554
rect 10089 6502 10141 6554
rect 10153 6502 10205 6554
rect 2780 6400 2832 6452
rect 3976 6400 4028 6452
rect 6092 6400 6144 6452
rect 3608 6332 3660 6384
rect 8116 6443 8168 6452
rect 8116 6409 8125 6443
rect 8125 6409 8159 6443
rect 8159 6409 8168 6443
rect 8116 6400 8168 6409
rect 9036 6400 9088 6452
rect 9864 6400 9916 6452
rect 10232 6400 10284 6452
rect 3516 6196 3568 6248
rect 5356 6264 5408 6316
rect 5632 6264 5684 6316
rect 8208 6332 8260 6384
rect 8392 6332 8444 6384
rect 7564 6307 7616 6316
rect 7564 6273 7573 6307
rect 7573 6273 7607 6307
rect 7607 6273 7616 6307
rect 7564 6264 7616 6273
rect 9496 6264 9548 6316
rect 5080 6196 5132 6248
rect 6828 6196 6880 6248
rect 8852 6239 8904 6248
rect 8852 6205 8861 6239
rect 8861 6205 8895 6239
rect 8895 6205 8904 6239
rect 8852 6196 8904 6205
rect 9128 6239 9180 6248
rect 9128 6205 9137 6239
rect 9137 6205 9171 6239
rect 9171 6205 9180 6239
rect 9128 6196 9180 6205
rect 4160 6128 4212 6180
rect 9680 6196 9732 6248
rect 10324 6128 10376 6180
rect 10784 6128 10836 6180
rect 2964 6060 3016 6112
rect 7932 6060 7984 6112
rect 9496 6060 9548 6112
rect 3112 5958 3164 6010
rect 3176 5958 3228 6010
rect 3240 5958 3292 6010
rect 3304 5958 3356 6010
rect 3368 5958 3420 6010
rect 5826 5958 5878 6010
rect 5890 5958 5942 6010
rect 5954 5958 6006 6010
rect 6018 5958 6070 6010
rect 6082 5958 6134 6010
rect 8540 5958 8592 6010
rect 8604 5958 8656 6010
rect 8668 5958 8720 6010
rect 8732 5958 8784 6010
rect 8796 5958 8848 6010
rect 11254 5958 11306 6010
rect 11318 5958 11370 6010
rect 11382 5958 11434 6010
rect 11446 5958 11498 6010
rect 11510 5958 11562 6010
rect 7656 5899 7708 5908
rect 7656 5865 7665 5899
rect 7665 5865 7699 5899
rect 7699 5865 7708 5899
rect 7656 5856 7708 5865
rect 9128 5856 9180 5908
rect 9220 5899 9272 5908
rect 9220 5865 9229 5899
rect 9229 5865 9263 5899
rect 9263 5865 9272 5899
rect 9220 5856 9272 5865
rect 10876 5856 10928 5908
rect 7564 5788 7616 5840
rect 8300 5788 8352 5840
rect 7748 5720 7800 5772
rect 8392 5720 8444 5772
rect 10232 5788 10284 5840
rect 8944 5720 8996 5772
rect 9496 5720 9548 5772
rect 9864 5763 9916 5772
rect 9864 5729 9873 5763
rect 9873 5729 9907 5763
rect 9907 5729 9916 5763
rect 9864 5720 9916 5729
rect 10600 5652 10652 5704
rect 9404 5627 9456 5636
rect 9404 5593 9413 5627
rect 9413 5593 9447 5627
rect 9447 5593 9456 5627
rect 9404 5584 9456 5593
rect 10508 5627 10560 5636
rect 10508 5593 10517 5627
rect 10517 5593 10551 5627
rect 10551 5593 10560 5627
rect 10508 5584 10560 5593
rect 1755 5414 1807 5466
rect 1819 5414 1871 5466
rect 1883 5414 1935 5466
rect 1947 5414 1999 5466
rect 2011 5414 2063 5466
rect 4469 5414 4521 5466
rect 4533 5414 4585 5466
rect 4597 5414 4649 5466
rect 4661 5414 4713 5466
rect 4725 5414 4777 5466
rect 7183 5414 7235 5466
rect 7247 5414 7299 5466
rect 7311 5414 7363 5466
rect 7375 5414 7427 5466
rect 7439 5414 7491 5466
rect 9897 5414 9949 5466
rect 9961 5414 10013 5466
rect 10025 5414 10077 5466
rect 10089 5414 10141 5466
rect 10153 5414 10205 5466
rect 10324 5355 10376 5364
rect 10324 5321 10333 5355
rect 10333 5321 10367 5355
rect 10367 5321 10376 5355
rect 10324 5312 10376 5321
rect 10600 5355 10652 5364
rect 10600 5321 10609 5355
rect 10609 5321 10643 5355
rect 10643 5321 10652 5355
rect 10600 5312 10652 5321
rect 10232 5244 10284 5296
rect 10416 5108 10468 5160
rect 10968 5040 11020 5092
rect 3112 4870 3164 4922
rect 3176 4870 3228 4922
rect 3240 4870 3292 4922
rect 3304 4870 3356 4922
rect 3368 4870 3420 4922
rect 5826 4870 5878 4922
rect 5890 4870 5942 4922
rect 5954 4870 6006 4922
rect 6018 4870 6070 4922
rect 6082 4870 6134 4922
rect 8540 4870 8592 4922
rect 8604 4870 8656 4922
rect 8668 4870 8720 4922
rect 8732 4870 8784 4922
rect 8796 4870 8848 4922
rect 11254 4870 11306 4922
rect 11318 4870 11370 4922
rect 11382 4870 11434 4922
rect 11446 4870 11498 4922
rect 11510 4870 11562 4922
rect 10784 4811 10836 4820
rect 10784 4777 10793 4811
rect 10793 4777 10827 4811
rect 10827 4777 10836 4811
rect 10784 4768 10836 4777
rect 10324 4700 10376 4752
rect 9496 4632 9548 4684
rect 10692 4675 10744 4684
rect 10692 4641 10701 4675
rect 10701 4641 10735 4675
rect 10735 4641 10744 4675
rect 10692 4632 10744 4641
rect 1755 4326 1807 4378
rect 1819 4326 1871 4378
rect 1883 4326 1935 4378
rect 1947 4326 1999 4378
rect 2011 4326 2063 4378
rect 4469 4326 4521 4378
rect 4533 4326 4585 4378
rect 4597 4326 4649 4378
rect 4661 4326 4713 4378
rect 4725 4326 4777 4378
rect 7183 4326 7235 4378
rect 7247 4326 7299 4378
rect 7311 4326 7363 4378
rect 7375 4326 7427 4378
rect 7439 4326 7491 4378
rect 9897 4326 9949 4378
rect 9961 4326 10013 4378
rect 10025 4326 10077 4378
rect 10089 4326 10141 4378
rect 10153 4326 10205 4378
rect 3112 3782 3164 3834
rect 3176 3782 3228 3834
rect 3240 3782 3292 3834
rect 3304 3782 3356 3834
rect 3368 3782 3420 3834
rect 5826 3782 5878 3834
rect 5890 3782 5942 3834
rect 5954 3782 6006 3834
rect 6018 3782 6070 3834
rect 6082 3782 6134 3834
rect 8540 3782 8592 3834
rect 8604 3782 8656 3834
rect 8668 3782 8720 3834
rect 8732 3782 8784 3834
rect 8796 3782 8848 3834
rect 11254 3782 11306 3834
rect 11318 3782 11370 3834
rect 11382 3782 11434 3834
rect 11446 3782 11498 3834
rect 11510 3782 11562 3834
rect 1755 3238 1807 3290
rect 1819 3238 1871 3290
rect 1883 3238 1935 3290
rect 1947 3238 1999 3290
rect 2011 3238 2063 3290
rect 4469 3238 4521 3290
rect 4533 3238 4585 3290
rect 4597 3238 4649 3290
rect 4661 3238 4713 3290
rect 4725 3238 4777 3290
rect 7183 3238 7235 3290
rect 7247 3238 7299 3290
rect 7311 3238 7363 3290
rect 7375 3238 7427 3290
rect 7439 3238 7491 3290
rect 9897 3238 9949 3290
rect 9961 3238 10013 3290
rect 10025 3238 10077 3290
rect 10089 3238 10141 3290
rect 10153 3238 10205 3290
rect 3112 2694 3164 2746
rect 3176 2694 3228 2746
rect 3240 2694 3292 2746
rect 3304 2694 3356 2746
rect 3368 2694 3420 2746
rect 5826 2694 5878 2746
rect 5890 2694 5942 2746
rect 5954 2694 6006 2746
rect 6018 2694 6070 2746
rect 6082 2694 6134 2746
rect 8540 2694 8592 2746
rect 8604 2694 8656 2746
rect 8668 2694 8720 2746
rect 8732 2694 8784 2746
rect 8796 2694 8848 2746
rect 11254 2694 11306 2746
rect 11318 2694 11370 2746
rect 11382 2694 11434 2746
rect 11446 2694 11498 2746
rect 11510 2694 11562 2746
rect 1755 2150 1807 2202
rect 1819 2150 1871 2202
rect 1883 2150 1935 2202
rect 1947 2150 1999 2202
rect 2011 2150 2063 2202
rect 4469 2150 4521 2202
rect 4533 2150 4585 2202
rect 4597 2150 4649 2202
rect 4661 2150 4713 2202
rect 4725 2150 4777 2202
rect 7183 2150 7235 2202
rect 7247 2150 7299 2202
rect 7311 2150 7363 2202
rect 7375 2150 7427 2202
rect 7439 2150 7491 2202
rect 9897 2150 9949 2202
rect 9961 2150 10013 2202
rect 10025 2150 10077 2202
rect 10089 2150 10141 2202
rect 10153 2150 10205 2202
rect 3112 1606 3164 1658
rect 3176 1606 3228 1658
rect 3240 1606 3292 1658
rect 3304 1606 3356 1658
rect 3368 1606 3420 1658
rect 5826 1606 5878 1658
rect 5890 1606 5942 1658
rect 5954 1606 6006 1658
rect 6018 1606 6070 1658
rect 6082 1606 6134 1658
rect 8540 1606 8592 1658
rect 8604 1606 8656 1658
rect 8668 1606 8720 1658
rect 8732 1606 8784 1658
rect 8796 1606 8848 1658
rect 11254 1606 11306 1658
rect 11318 1606 11370 1658
rect 11382 1606 11434 1658
rect 11446 1606 11498 1658
rect 11510 1606 11562 1658
rect 1755 1062 1807 1114
rect 1819 1062 1871 1114
rect 1883 1062 1935 1114
rect 1947 1062 1999 1114
rect 2011 1062 2063 1114
rect 4469 1062 4521 1114
rect 4533 1062 4585 1114
rect 4597 1062 4649 1114
rect 4661 1062 4713 1114
rect 4725 1062 4777 1114
rect 7183 1062 7235 1114
rect 7247 1062 7299 1114
rect 7311 1062 7363 1114
rect 7375 1062 7427 1114
rect 7439 1062 7491 1114
rect 9897 1062 9949 1114
rect 9961 1062 10013 1114
rect 10025 1062 10077 1114
rect 10089 1062 10141 1114
rect 10153 1062 10205 1114
rect 3112 518 3164 570
rect 3176 518 3228 570
rect 3240 518 3292 570
rect 3304 518 3356 570
rect 3368 518 3420 570
rect 5826 518 5878 570
rect 5890 518 5942 570
rect 5954 518 6006 570
rect 6018 518 6070 570
rect 6082 518 6134 570
rect 8540 518 8592 570
rect 8604 518 8656 570
rect 8668 518 8720 570
rect 8732 518 8784 570
rect 8796 518 8848 570
rect 11254 518 11306 570
rect 11318 518 11370 570
rect 11382 518 11434 570
rect 11446 518 11498 570
rect 11510 518 11562 570
<< metal2 >>
rect 754 11600 810 12000
rect 2042 11600 2098 12000
rect 3330 11600 3386 12000
rect 3976 11688 4028 11694
rect 3976 11630 4028 11636
rect 768 10810 796 11600
rect 2056 11098 2084 11600
rect 3344 11558 3372 11600
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 3332 11552 3384 11558
rect 3332 11494 3384 11500
rect 2688 11280 2740 11286
rect 2688 11222 2740 11228
rect 2056 11070 2176 11098
rect 1755 10908 2063 10917
rect 1755 10906 1761 10908
rect 1817 10906 1841 10908
rect 1897 10906 1921 10908
rect 1977 10906 2001 10908
rect 2057 10906 2063 10908
rect 1817 10854 1819 10906
rect 1999 10854 2001 10906
rect 1755 10852 1761 10854
rect 1817 10852 1841 10854
rect 1897 10852 1921 10854
rect 1977 10852 2001 10854
rect 2057 10852 2063 10854
rect 1755 10843 2063 10852
rect 2148 10810 2176 11070
rect 756 10804 808 10810
rect 756 10746 808 10752
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 1032 10736 1084 10742
rect 1032 10678 1084 10684
rect 1044 10130 1072 10678
rect 1308 10600 1360 10606
rect 1308 10542 1360 10548
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1216 10532 1268 10538
rect 1216 10474 1268 10480
rect 1124 10192 1176 10198
rect 1124 10134 1176 10140
rect 1032 10124 1084 10130
rect 1032 10066 1084 10072
rect 1136 9654 1164 10134
rect 1228 10130 1256 10474
rect 1216 10124 1268 10130
rect 1216 10066 1268 10072
rect 1216 9920 1268 9926
rect 1216 9862 1268 9868
rect 1124 9648 1176 9654
rect 1228 9625 1256 9862
rect 1320 9722 1348 10542
rect 1688 9994 1716 10542
rect 2596 10464 2648 10470
rect 2596 10406 2648 10412
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 1676 9988 1728 9994
rect 1676 9930 1728 9936
rect 1584 9920 1636 9926
rect 1584 9862 1636 9868
rect 1308 9716 1360 9722
rect 1308 9658 1360 9664
rect 1124 9590 1176 9596
rect 1214 9616 1270 9625
rect 1214 9551 1270 9560
rect 1596 9518 1624 9862
rect 1755 9820 2063 9829
rect 1755 9818 1761 9820
rect 1817 9818 1841 9820
rect 1897 9818 1921 9820
rect 1977 9818 2001 9820
rect 2057 9818 2063 9820
rect 1817 9766 1819 9818
rect 1999 9766 2001 9818
rect 1755 9764 1761 9766
rect 1817 9764 1841 9766
rect 1897 9764 1921 9766
rect 1977 9764 2001 9766
rect 2057 9764 2063 9766
rect 1755 9755 2063 9764
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 2424 9178 2452 10066
rect 2608 9382 2636 10406
rect 2700 10266 2728 11222
rect 2884 10810 2912 11494
rect 3112 11452 3420 11461
rect 3112 11450 3118 11452
rect 3174 11450 3198 11452
rect 3254 11450 3278 11452
rect 3334 11450 3358 11452
rect 3414 11450 3420 11452
rect 3174 11398 3176 11450
rect 3356 11398 3358 11450
rect 3112 11396 3118 11398
rect 3174 11396 3198 11398
rect 3254 11396 3278 11398
rect 3334 11396 3358 11398
rect 3414 11396 3420 11398
rect 3112 11387 3420 11396
rect 3988 11286 4016 11630
rect 4618 11600 4674 12000
rect 5906 11600 5962 12000
rect 6644 11620 6696 11626
rect 4632 11354 4660 11600
rect 5920 11558 5948 11600
rect 7194 11600 7250 12000
rect 7840 11688 7892 11694
rect 7840 11630 7892 11636
rect 6644 11562 6696 11568
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 5826 11452 6134 11461
rect 5826 11450 5832 11452
rect 5888 11450 5912 11452
rect 5968 11450 5992 11452
rect 6048 11450 6072 11452
rect 6128 11450 6134 11452
rect 5888 11398 5890 11450
rect 6070 11398 6072 11450
rect 5826 11396 5832 11398
rect 5888 11396 5912 11398
rect 5968 11396 5992 11398
rect 6048 11396 6072 11398
rect 6128 11396 6134 11398
rect 5826 11387 6134 11396
rect 6196 11354 6224 11494
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 3976 11280 4028 11286
rect 3976 11222 4028 11228
rect 3056 11212 3108 11218
rect 3056 11154 3108 11160
rect 2964 11008 3016 11014
rect 2964 10950 3016 10956
rect 2872 10804 2924 10810
rect 2872 10746 2924 10752
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2872 10192 2924 10198
rect 2872 10134 2924 10140
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2608 8906 2636 9318
rect 2596 8900 2648 8906
rect 2596 8842 2648 8848
rect 1755 8732 2063 8741
rect 1755 8730 1761 8732
rect 1817 8730 1841 8732
rect 1897 8730 1921 8732
rect 1977 8730 2001 8732
rect 2057 8730 2063 8732
rect 1817 8678 1819 8730
rect 1999 8678 2001 8730
rect 1755 8676 1761 8678
rect 1817 8676 1841 8678
rect 1897 8676 1921 8678
rect 1977 8676 2001 8678
rect 2057 8676 2063 8678
rect 1755 8667 2063 8676
rect 2792 8634 2820 10066
rect 2884 9178 2912 10134
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 2976 8430 3004 10950
rect 3068 10810 3096 11154
rect 3608 11144 3660 11150
rect 3608 11086 3660 11092
rect 3792 11144 3844 11150
rect 3792 11086 3844 11092
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 3068 10606 3096 10746
rect 3620 10606 3648 11086
rect 3700 11008 3752 11014
rect 3700 10950 3752 10956
rect 3712 10606 3740 10950
rect 3804 10742 3832 11086
rect 3988 10826 4016 11222
rect 6656 11218 6684 11562
rect 7208 11558 7236 11600
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 7024 11342 7236 11370
rect 7024 11234 7052 11342
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6840 11206 7052 11234
rect 7104 11212 7156 11218
rect 4988 11008 5040 11014
rect 4988 10950 5040 10956
rect 4469 10908 4777 10917
rect 4469 10906 4475 10908
rect 4531 10906 4555 10908
rect 4611 10906 4635 10908
rect 4691 10906 4715 10908
rect 4771 10906 4777 10908
rect 4531 10854 4533 10906
rect 4713 10854 4715 10906
rect 4469 10852 4475 10854
rect 4531 10852 4555 10854
rect 4611 10852 4635 10854
rect 4691 10852 4715 10854
rect 4771 10852 4777 10854
rect 4469 10843 4777 10852
rect 3988 10798 4200 10826
rect 3792 10736 3844 10742
rect 3792 10678 3844 10684
rect 4068 10736 4120 10742
rect 4068 10678 4120 10684
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 3240 10600 3292 10606
rect 3240 10542 3292 10548
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 3700 10600 3752 10606
rect 3700 10542 3752 10548
rect 3252 10452 3280 10542
rect 3252 10424 3556 10452
rect 3112 10364 3420 10373
rect 3112 10362 3118 10364
rect 3174 10362 3198 10364
rect 3254 10362 3278 10364
rect 3334 10362 3358 10364
rect 3414 10362 3420 10364
rect 3174 10310 3176 10362
rect 3356 10310 3358 10362
rect 3112 10308 3118 10310
rect 3174 10308 3198 10310
rect 3254 10308 3278 10310
rect 3334 10308 3358 10310
rect 3414 10308 3420 10310
rect 3112 10299 3420 10308
rect 3528 10266 3556 10424
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 3424 10124 3476 10130
rect 3424 10066 3476 10072
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 3068 9654 3096 9998
rect 3056 9648 3108 9654
rect 3056 9590 3108 9596
rect 3330 9616 3386 9625
rect 3330 9551 3386 9560
rect 3056 9512 3108 9518
rect 3054 9480 3056 9489
rect 3108 9480 3110 9489
rect 3344 9450 3372 9551
rect 3054 9415 3110 9424
rect 3332 9444 3384 9450
rect 3436 9432 3464 10066
rect 3620 9926 3648 10542
rect 3712 10266 3740 10542
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3516 9512 3568 9518
rect 3568 9460 3740 9466
rect 3516 9454 3740 9460
rect 3528 9438 3740 9454
rect 3436 9404 3496 9432
rect 3332 9386 3384 9392
rect 3468 9364 3496 9404
rect 3468 9336 3556 9364
rect 3112 9276 3420 9285
rect 3112 9274 3118 9276
rect 3174 9274 3198 9276
rect 3254 9274 3278 9276
rect 3334 9274 3358 9276
rect 3414 9274 3420 9276
rect 3174 9222 3176 9274
rect 3356 9222 3358 9274
rect 3112 9220 3118 9222
rect 3174 9220 3198 9222
rect 3254 9220 3278 9222
rect 3334 9220 3358 9222
rect 3414 9220 3420 9222
rect 3112 9211 3420 9220
rect 3332 8832 3384 8838
rect 3528 8820 3556 9336
rect 3712 8974 3740 9438
rect 3804 9178 3832 10678
rect 3976 10600 4028 10606
rect 3976 10542 4028 10548
rect 3884 9920 3936 9926
rect 3988 9874 4016 10542
rect 3936 9868 4016 9874
rect 3884 9862 4016 9868
rect 3896 9846 4016 9862
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 3988 9110 4016 9846
rect 4080 9382 4108 10678
rect 4172 10606 4200 10798
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 4172 10130 4200 10542
rect 4804 10532 4856 10538
rect 4804 10474 4856 10480
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 3976 9104 4028 9110
rect 3976 9046 4028 9052
rect 3700 8968 3752 8974
rect 3700 8910 3752 8916
rect 3384 8792 3556 8820
rect 3332 8774 3384 8780
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 3344 8362 3372 8774
rect 3516 8560 3568 8566
rect 3516 8502 3568 8508
rect 3332 8356 3384 8362
rect 3332 8298 3384 8304
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2976 7954 3004 8230
rect 3112 8188 3420 8197
rect 3112 8186 3118 8188
rect 3174 8186 3198 8188
rect 3254 8186 3278 8188
rect 3334 8186 3358 8188
rect 3414 8186 3420 8188
rect 3174 8134 3176 8186
rect 3356 8134 3358 8186
rect 3112 8132 3118 8134
rect 3174 8132 3198 8134
rect 3254 8132 3278 8134
rect 3334 8132 3358 8134
rect 3414 8132 3420 8134
rect 3112 8123 3420 8132
rect 3528 7970 3556 8502
rect 3608 8424 3660 8430
rect 3608 8366 3660 8372
rect 3436 7954 3556 7970
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 3424 7948 3556 7954
rect 3476 7942 3556 7948
rect 3424 7890 3476 7896
rect 2596 7744 2648 7750
rect 2596 7686 2648 7692
rect 1755 7644 2063 7653
rect 1755 7642 1761 7644
rect 1817 7642 1841 7644
rect 1897 7642 1921 7644
rect 1977 7642 2001 7644
rect 2057 7642 2063 7644
rect 1817 7590 1819 7642
rect 1999 7590 2001 7642
rect 1755 7588 1761 7590
rect 1817 7588 1841 7590
rect 1897 7588 1921 7590
rect 1977 7588 2001 7590
rect 2057 7588 2063 7590
rect 1755 7579 2063 7588
rect 2608 7410 2636 7686
rect 2596 7404 2648 7410
rect 2596 7346 2648 7352
rect 2504 7268 2556 7274
rect 2504 7210 2556 7216
rect 2516 6866 2544 7210
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 1755 6556 2063 6565
rect 1755 6554 1761 6556
rect 1817 6554 1841 6556
rect 1897 6554 1921 6556
rect 1977 6554 2001 6556
rect 2057 6554 2063 6556
rect 1817 6502 1819 6554
rect 1999 6502 2001 6554
rect 1755 6500 1761 6502
rect 1817 6500 1841 6502
rect 1897 6500 1921 6502
rect 1977 6500 2001 6502
rect 2057 6500 2063 6502
rect 1755 6491 2063 6500
rect 2792 6458 2820 7890
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 2976 7546 3004 7686
rect 2964 7540 3016 7546
rect 2964 7482 3016 7488
rect 3344 7274 3372 7686
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 2964 7268 3016 7274
rect 2964 7210 3016 7216
rect 3332 7268 3384 7274
rect 3332 7210 3384 7216
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 2976 6118 3004 7210
rect 3112 7100 3420 7109
rect 3112 7098 3118 7100
rect 3174 7098 3198 7100
rect 3254 7098 3278 7100
rect 3334 7098 3358 7100
rect 3414 7098 3420 7100
rect 3174 7046 3176 7098
rect 3356 7046 3358 7098
rect 3112 7044 3118 7046
rect 3174 7044 3198 7046
rect 3254 7044 3278 7046
rect 3334 7044 3358 7046
rect 3414 7044 3420 7046
rect 3112 7035 3420 7044
rect 3528 7002 3556 7482
rect 3620 7206 3648 8366
rect 3712 8022 3740 8910
rect 3988 8430 4016 9046
rect 4080 8838 4108 9318
rect 4172 9042 4200 10066
rect 4816 10062 4844 10474
rect 5000 10198 5028 10950
rect 4988 10192 5040 10198
rect 4988 10134 5040 10140
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4469 9820 4777 9829
rect 4469 9818 4475 9820
rect 4531 9818 4555 9820
rect 4611 9818 4635 9820
rect 4691 9818 4715 9820
rect 4771 9818 4777 9820
rect 4531 9766 4533 9818
rect 4713 9766 4715 9818
rect 4469 9764 4475 9766
rect 4531 9764 4555 9766
rect 4611 9764 4635 9766
rect 4691 9764 4715 9766
rect 4771 9764 4777 9766
rect 4469 9755 4777 9764
rect 4816 9586 4844 9998
rect 4896 9648 4948 9654
rect 4896 9590 4948 9596
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 4908 9450 4936 9590
rect 4896 9444 4948 9450
rect 4896 9386 4948 9392
rect 4160 9036 4212 9042
rect 4212 8996 4292 9024
rect 4160 8978 4212 8984
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 4068 8560 4120 8566
rect 4120 8520 4200 8548
rect 4068 8502 4120 8508
rect 3976 8424 4028 8430
rect 3976 8366 4028 8372
rect 4172 8362 4200 8520
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 3700 8016 3752 8022
rect 3700 7958 3752 7964
rect 3712 7342 3740 7958
rect 3804 7342 3832 8230
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 3608 7200 3660 7206
rect 3608 7142 3660 7148
rect 3516 6996 3568 7002
rect 3516 6938 3568 6944
rect 3528 6254 3556 6938
rect 3620 6390 3648 7142
rect 3712 6798 3740 7278
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 3700 6792 3752 6798
rect 3700 6734 3752 6740
rect 3988 6458 4016 6802
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 3608 6384 3660 6390
rect 3608 6326 3660 6332
rect 3516 6248 3568 6254
rect 3516 6190 3568 6196
rect 4172 6186 4200 8298
rect 4264 6866 4292 8996
rect 4469 8732 4777 8741
rect 4469 8730 4475 8732
rect 4531 8730 4555 8732
rect 4611 8730 4635 8732
rect 4691 8730 4715 8732
rect 4771 8730 4777 8732
rect 4531 8678 4533 8730
rect 4713 8678 4715 8730
rect 4469 8676 4475 8678
rect 4531 8676 4555 8678
rect 4611 8676 4635 8678
rect 4691 8676 4715 8678
rect 4771 8676 4777 8678
rect 4469 8667 4777 8676
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4724 8090 4752 8434
rect 4804 8356 4856 8362
rect 4908 8344 4936 9386
rect 5184 8566 5212 11154
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5356 10532 5408 10538
rect 5356 10474 5408 10480
rect 5368 10266 5396 10474
rect 5356 10260 5408 10266
rect 5356 10202 5408 10208
rect 5552 10130 5580 11018
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 6748 10810 6776 10950
rect 6736 10804 6788 10810
rect 6736 10746 6788 10752
rect 6840 10554 6868 11206
rect 7104 11154 7156 11160
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 6932 10742 6960 11086
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 5724 10532 5776 10538
rect 6840 10526 6960 10554
rect 5724 10474 5776 10480
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5446 10024 5502 10033
rect 5446 9959 5502 9968
rect 5460 9654 5488 9959
rect 5448 9648 5500 9654
rect 5448 9590 5500 9596
rect 5448 9512 5500 9518
rect 5262 9480 5318 9489
rect 5448 9454 5500 9460
rect 5262 9415 5264 9424
rect 5316 9415 5318 9424
rect 5264 9386 5316 9392
rect 5460 8974 5488 9454
rect 5736 9178 5764 10474
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 5826 10364 6134 10373
rect 5826 10362 5832 10364
rect 5888 10362 5912 10364
rect 5968 10362 5992 10364
rect 6048 10362 6072 10364
rect 6128 10362 6134 10364
rect 5888 10310 5890 10362
rect 6070 10310 6072 10362
rect 5826 10308 5832 10310
rect 5888 10308 5912 10310
rect 5968 10308 5992 10310
rect 6048 10308 6072 10310
rect 6128 10308 6134 10310
rect 5826 10299 6134 10308
rect 6748 10198 6776 10406
rect 6736 10192 6788 10198
rect 6736 10134 6788 10140
rect 5816 9920 5868 9926
rect 5816 9862 5868 9868
rect 5828 9674 5856 9862
rect 6932 9674 6960 10526
rect 7024 10130 7052 11086
rect 7116 10470 7144 11154
rect 7208 11150 7236 11342
rect 7656 11280 7708 11286
rect 7708 11240 7788 11268
rect 7656 11222 7708 11228
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7196 11144 7248 11150
rect 7576 11098 7604 11154
rect 7196 11086 7248 11092
rect 7300 11082 7604 11098
rect 7288 11076 7604 11082
rect 7340 11070 7604 11076
rect 7656 11076 7708 11082
rect 7288 11018 7340 11024
rect 7656 11018 7708 11024
rect 7564 11008 7616 11014
rect 7564 10950 7616 10956
rect 7183 10908 7491 10917
rect 7183 10906 7189 10908
rect 7245 10906 7269 10908
rect 7325 10906 7349 10908
rect 7405 10906 7429 10908
rect 7485 10906 7491 10908
rect 7245 10854 7247 10906
rect 7427 10854 7429 10906
rect 7183 10852 7189 10854
rect 7245 10852 7269 10854
rect 7325 10852 7349 10854
rect 7405 10852 7429 10854
rect 7485 10852 7491 10854
rect 7183 10843 7491 10852
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 7024 9926 7052 10066
rect 7116 9994 7144 10406
rect 7484 10146 7512 10542
rect 7576 10266 7604 10950
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7484 10118 7604 10146
rect 7668 10130 7696 11018
rect 7760 11014 7788 11240
rect 7852 11218 7880 11630
rect 8024 11620 8076 11626
rect 8024 11562 8076 11568
rect 8300 11620 8352 11626
rect 8482 11620 8538 12000
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 8482 11600 8484 11620
rect 8300 11562 8352 11568
rect 8536 11600 8538 11620
rect 8484 11562 8536 11568
rect 8036 11218 8064 11562
rect 8312 11354 8340 11562
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 8540 11452 8848 11461
rect 8540 11450 8546 11452
rect 8602 11450 8626 11452
rect 8682 11450 8706 11452
rect 8762 11450 8786 11452
rect 8842 11450 8848 11452
rect 8602 11398 8604 11450
rect 8784 11398 8786 11450
rect 8540 11396 8546 11398
rect 8602 11396 8626 11398
rect 8682 11396 8706 11398
rect 8762 11396 8786 11398
rect 8842 11396 8848 11398
rect 8540 11387 8848 11396
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 7840 11212 7892 11218
rect 7840 11154 7892 11160
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 7932 11076 7984 11082
rect 7932 11018 7984 11024
rect 7748 11008 7800 11014
rect 7748 10950 7800 10956
rect 7760 10606 7788 10950
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 7024 9722 7052 9862
rect 7183 9820 7491 9829
rect 7183 9818 7189 9820
rect 7245 9818 7269 9820
rect 7325 9818 7349 9820
rect 7405 9818 7429 9820
rect 7485 9818 7491 9820
rect 7245 9766 7247 9818
rect 7427 9766 7429 9818
rect 7183 9764 7189 9766
rect 7245 9764 7269 9766
rect 7325 9764 7349 9766
rect 7405 9764 7429 9766
rect 7485 9764 7491 9766
rect 7183 9755 7491 9764
rect 5828 9646 5948 9674
rect 5920 9450 5948 9646
rect 6840 9646 6960 9674
rect 7012 9716 7064 9722
rect 7012 9658 7064 9664
rect 7288 9648 7340 9654
rect 6840 9489 6868 9646
rect 7288 9590 7340 9596
rect 7300 9489 7328 9590
rect 6826 9480 6882 9489
rect 5908 9444 5960 9450
rect 6826 9415 6882 9424
rect 7286 9480 7342 9489
rect 7576 9450 7604 10118
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7760 10010 7788 10542
rect 7944 10470 7972 11018
rect 8036 10674 8064 11154
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 7668 9982 7788 10010
rect 7286 9415 7342 9424
rect 7564 9444 7616 9450
rect 5908 9386 5960 9392
rect 5826 9276 6134 9285
rect 5826 9274 5832 9276
rect 5888 9274 5912 9276
rect 5968 9274 5992 9276
rect 6048 9274 6072 9276
rect 6128 9274 6134 9276
rect 5888 9222 5890 9274
rect 6070 9222 6072 9274
rect 5826 9220 5832 9222
rect 5888 9220 5912 9222
rect 5968 9220 5992 9222
rect 6048 9220 6072 9222
rect 6128 9220 6134 9222
rect 5826 9211 6134 9220
rect 5724 9172 5776 9178
rect 5724 9114 5776 9120
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5172 8560 5224 8566
rect 5172 8502 5224 8508
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 6276 8424 6328 8430
rect 6276 8366 6328 8372
rect 4856 8316 4936 8344
rect 4988 8356 5040 8362
rect 4804 8298 4856 8304
rect 4988 8298 5040 8304
rect 5080 8356 5132 8362
rect 5080 8298 5132 8304
rect 4712 8084 4764 8090
rect 4712 8026 4764 8032
rect 5000 7750 5028 8298
rect 4988 7744 5040 7750
rect 4988 7686 5040 7692
rect 4469 7644 4777 7653
rect 4469 7642 4475 7644
rect 4531 7642 4555 7644
rect 4611 7642 4635 7644
rect 4691 7642 4715 7644
rect 4771 7642 4777 7644
rect 4531 7590 4533 7642
rect 4713 7590 4715 7642
rect 4469 7588 4475 7590
rect 4531 7588 4555 7590
rect 4611 7588 4635 7590
rect 4691 7588 4715 7590
rect 4771 7588 4777 7590
rect 4469 7579 4777 7588
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 5092 6730 5120 8298
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5184 7546 5212 8230
rect 5276 7954 5304 8230
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5184 7342 5212 7482
rect 5276 7342 5304 7890
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5368 7206 5396 7686
rect 5460 7546 5488 7822
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5552 7342 5580 7686
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 5644 6934 5672 7278
rect 5632 6928 5684 6934
rect 5632 6870 5684 6876
rect 5080 6724 5132 6730
rect 5080 6666 5132 6672
rect 4469 6556 4777 6565
rect 4469 6554 4475 6556
rect 4531 6554 4555 6556
rect 4611 6554 4635 6556
rect 4691 6554 4715 6556
rect 4771 6554 4777 6556
rect 4531 6502 4533 6554
rect 4713 6502 4715 6554
rect 4469 6500 4475 6502
rect 4531 6500 4555 6502
rect 4611 6500 4635 6502
rect 4691 6500 4715 6502
rect 4771 6500 4777 6502
rect 4469 6491 4777 6500
rect 5092 6254 5120 6666
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5368 6322 5396 6598
rect 5644 6322 5672 6870
rect 5736 6866 5764 8366
rect 6184 8288 6236 8294
rect 6184 8230 6236 8236
rect 5826 8188 6134 8197
rect 5826 8186 5832 8188
rect 5888 8186 5912 8188
rect 5968 8186 5992 8188
rect 6048 8186 6072 8188
rect 6128 8186 6134 8188
rect 5888 8134 5890 8186
rect 6070 8134 6072 8186
rect 5826 8132 5832 8134
rect 5888 8132 5912 8134
rect 5968 8132 5992 8134
rect 6048 8132 6072 8134
rect 6128 8132 6134 8134
rect 5826 8123 6134 8132
rect 6196 7342 6224 8230
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 5826 7100 6134 7109
rect 5826 7098 5832 7100
rect 5888 7098 5912 7100
rect 5968 7098 5992 7100
rect 6048 7098 6072 7100
rect 6128 7098 6134 7100
rect 5888 7046 5890 7098
rect 6070 7046 6072 7098
rect 5826 7044 5832 7046
rect 5888 7044 5912 7046
rect 5968 7044 5992 7046
rect 6048 7044 6072 7046
rect 6128 7044 6134 7046
rect 5826 7035 6134 7044
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 6104 6458 6132 6802
rect 6288 6730 6316 8366
rect 6380 7750 6408 8978
rect 6840 8430 6868 9415
rect 7564 9386 7616 9392
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7288 9376 7340 9382
rect 7668 9330 7696 9982
rect 7748 9920 7800 9926
rect 7852 9874 7880 10066
rect 7800 9868 7880 9874
rect 7748 9862 7880 9868
rect 7760 9846 7880 9862
rect 7760 9586 7788 9846
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7340 9324 7696 9330
rect 7288 9318 7696 9324
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 6460 8424 6512 8430
rect 6828 8424 6880 8430
rect 6460 8366 6512 8372
rect 6748 8384 6828 8412
rect 6472 8090 6500 8366
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6656 6866 6684 8298
rect 6748 7274 6776 8384
rect 6828 8366 6880 8372
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6736 7268 6788 7274
rect 6736 7210 6788 7216
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6276 6724 6328 6730
rect 6276 6666 6328 6672
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 6840 6254 6868 8230
rect 6932 8090 6960 8366
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 7024 7426 7052 8570
rect 7116 8498 7144 9318
rect 7300 9302 7696 9318
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7183 8732 7491 8741
rect 7183 8730 7189 8732
rect 7245 8730 7269 8732
rect 7325 8730 7349 8732
rect 7405 8730 7429 8732
rect 7485 8730 7491 8732
rect 7245 8678 7247 8730
rect 7427 8678 7429 8730
rect 7183 8676 7189 8678
rect 7245 8676 7269 8678
rect 7325 8676 7349 8678
rect 7405 8676 7429 8678
rect 7485 8676 7491 8678
rect 7183 8667 7491 8676
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7208 7886 7236 8366
rect 7484 8106 7512 8366
rect 7668 8106 7696 8774
rect 7760 8634 7788 9318
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7760 8430 7788 8570
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 7484 8090 7604 8106
rect 7484 8084 7616 8090
rect 7484 8078 7564 8084
rect 7484 7886 7512 8078
rect 7668 8078 7788 8106
rect 7564 8026 7616 8032
rect 7656 8016 7708 8022
rect 7656 7958 7708 7964
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7208 7732 7236 7822
rect 7116 7704 7236 7732
rect 7116 7546 7144 7704
rect 7183 7644 7491 7653
rect 7183 7642 7189 7644
rect 7245 7642 7269 7644
rect 7325 7642 7349 7644
rect 7405 7642 7429 7644
rect 7485 7642 7491 7644
rect 7245 7590 7247 7642
rect 7427 7590 7429 7642
rect 7183 7588 7189 7590
rect 7245 7588 7269 7590
rect 7325 7588 7349 7590
rect 7405 7588 7429 7590
rect 7485 7588 7491 7590
rect 7183 7579 7491 7588
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 7024 7398 7144 7426
rect 7116 7342 7144 7398
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 7116 6934 7144 7278
rect 7104 6928 7156 6934
rect 7104 6870 7156 6876
rect 7183 6556 7491 6565
rect 7183 6554 7189 6556
rect 7245 6554 7269 6556
rect 7325 6554 7349 6556
rect 7405 6554 7429 6556
rect 7485 6554 7491 6556
rect 7245 6502 7247 6554
rect 7427 6502 7429 6554
rect 7183 6500 7189 6502
rect 7245 6500 7269 6502
rect 7325 6500 7349 6502
rect 7405 6500 7429 6502
rect 7485 6500 7491 6502
rect 7183 6491 7491 6500
rect 7576 6322 7604 7890
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 5080 6248 5132 6254
rect 5080 6190 5132 6196
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 4160 6180 4212 6186
rect 4160 6122 4212 6128
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 3112 6012 3420 6021
rect 3112 6010 3118 6012
rect 3174 6010 3198 6012
rect 3254 6010 3278 6012
rect 3334 6010 3358 6012
rect 3414 6010 3420 6012
rect 3174 5958 3176 6010
rect 3356 5958 3358 6010
rect 3112 5956 3118 5958
rect 3174 5956 3198 5958
rect 3254 5956 3278 5958
rect 3334 5956 3358 5958
rect 3414 5956 3420 5958
rect 3112 5947 3420 5956
rect 5826 6012 6134 6021
rect 5826 6010 5832 6012
rect 5888 6010 5912 6012
rect 5968 6010 5992 6012
rect 6048 6010 6072 6012
rect 6128 6010 6134 6012
rect 5888 5958 5890 6010
rect 6070 5958 6072 6010
rect 5826 5956 5832 5958
rect 5888 5956 5912 5958
rect 5968 5956 5992 5958
rect 6048 5956 6072 5958
rect 6128 5956 6134 5958
rect 5826 5947 6134 5956
rect 7576 5846 7604 6258
rect 7668 5914 7696 7958
rect 7760 7818 7788 8078
rect 7748 7812 7800 7818
rect 7748 7754 7800 7760
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 7760 6662 7788 7278
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7564 5840 7616 5846
rect 7564 5782 7616 5788
rect 7760 5778 7788 6598
rect 7852 5817 7880 8978
rect 7944 8974 7972 10406
rect 8036 9926 8064 10610
rect 8128 10266 8156 11086
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8208 10736 8260 10742
rect 8208 10678 8260 10684
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 8220 10130 8248 10678
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8312 9994 8340 10746
rect 8540 10364 8848 10373
rect 8540 10362 8546 10364
rect 8602 10362 8626 10364
rect 8682 10362 8706 10364
rect 8762 10362 8786 10364
rect 8842 10362 8848 10364
rect 8602 10310 8604 10362
rect 8784 10310 8786 10362
rect 8540 10308 8546 10310
rect 8602 10308 8626 10310
rect 8682 10308 8706 10310
rect 8762 10308 8786 10310
rect 8842 10308 8848 10310
rect 8540 10299 8848 10308
rect 8300 9988 8352 9994
rect 8300 9930 8352 9936
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 8116 9444 8168 9450
rect 8116 9386 8168 9392
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 7944 7546 7972 8366
rect 8036 8022 8064 9318
rect 8128 8838 8156 9386
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 8220 8650 8248 9658
rect 8312 9654 8340 9930
rect 8956 9722 8984 11154
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 8944 9716 8996 9722
rect 8944 9658 8996 9664
rect 8300 9648 8352 9654
rect 9324 9625 9352 10406
rect 9508 10266 9536 11494
rect 9600 10266 9628 11630
rect 9770 11600 9826 12000
rect 11058 11600 11114 12000
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9680 10192 9732 10198
rect 9680 10134 9732 10140
rect 8300 9590 8352 9596
rect 9310 9616 9366 9625
rect 9310 9551 9366 9560
rect 9692 9518 9720 10134
rect 9784 10033 9812 11600
rect 11072 11370 11100 11600
rect 11254 11452 11562 11461
rect 11254 11450 11260 11452
rect 11316 11450 11340 11452
rect 11396 11450 11420 11452
rect 11476 11450 11500 11452
rect 11556 11450 11562 11452
rect 11316 11398 11318 11450
rect 11498 11398 11500 11450
rect 11254 11396 11260 11398
rect 11316 11396 11340 11398
rect 11396 11396 11420 11398
rect 11476 11396 11500 11398
rect 11556 11396 11562 11398
rect 11254 11387 11562 11396
rect 11072 11342 11192 11370
rect 11060 11280 11112 11286
rect 11060 11222 11112 11228
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 9897 10908 10205 10917
rect 9897 10906 9903 10908
rect 9959 10906 9983 10908
rect 10039 10906 10063 10908
rect 10119 10906 10143 10908
rect 10199 10906 10205 10908
rect 9959 10854 9961 10906
rect 10141 10854 10143 10906
rect 9897 10852 9903 10854
rect 9959 10852 9983 10854
rect 10039 10852 10063 10854
rect 10119 10852 10143 10854
rect 10199 10852 10205 10854
rect 9897 10843 10205 10852
rect 9770 10024 9826 10033
rect 9770 9959 9826 9968
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 8668 9512 8720 9518
rect 8666 9480 8668 9489
rect 9680 9512 9732 9518
rect 8720 9480 8722 9489
rect 9680 9454 9732 9460
rect 8666 9415 8722 9424
rect 9036 9444 9088 9450
rect 9036 9386 9088 9392
rect 8540 9276 8848 9285
rect 8540 9274 8546 9276
rect 8602 9274 8626 9276
rect 8682 9274 8706 9276
rect 8762 9274 8786 9276
rect 8842 9274 8848 9276
rect 8602 9222 8604 9274
rect 8784 9222 8786 9274
rect 8540 9220 8546 9222
rect 8602 9220 8626 9222
rect 8682 9220 8706 9222
rect 8762 9220 8786 9222
rect 8842 9220 8848 9222
rect 8540 9211 8848 9220
rect 9048 9178 9076 9386
rect 9036 9172 9088 9178
rect 9036 9114 9088 9120
rect 9784 8974 9812 9862
rect 9897 9820 10205 9829
rect 9897 9818 9903 9820
rect 9959 9818 9983 9820
rect 10039 9818 10063 9820
rect 10119 9818 10143 9820
rect 10199 9818 10205 9820
rect 9959 9766 9961 9818
rect 10141 9766 10143 9818
rect 9897 9764 9903 9766
rect 9959 9764 9983 9766
rect 10039 9764 10063 9766
rect 10119 9764 10143 9766
rect 10199 9764 10205 9766
rect 9897 9755 10205 9764
rect 10244 9382 10272 10950
rect 10796 10674 10824 11086
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 11072 10606 11100 11222
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10324 9512 10376 9518
rect 10324 9454 10376 9460
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 10336 9110 10364 9454
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10324 9104 10376 9110
rect 10324 9046 10376 9052
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8128 8622 8248 8650
rect 8128 8090 8156 8622
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 8116 8084 8168 8090
rect 8116 8026 8168 8032
rect 8024 8016 8076 8022
rect 8220 7970 8248 8366
rect 8024 7958 8076 7964
rect 8128 7942 8248 7970
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 7932 7268 7984 7274
rect 7932 7210 7984 7216
rect 7944 6118 7972 7210
rect 8128 7206 8156 7942
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8220 7546 8248 7822
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8208 7268 8260 7274
rect 8208 7210 8260 7216
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8128 6458 8156 7142
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8220 6390 8248 7210
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 8312 5846 8340 8774
rect 9897 8732 10205 8741
rect 9897 8730 9903 8732
rect 9959 8730 9983 8732
rect 10039 8730 10063 8732
rect 10119 8730 10143 8732
rect 10199 8730 10205 8732
rect 9959 8678 9961 8730
rect 10141 8678 10143 8730
rect 9897 8676 9903 8678
rect 9959 8676 9983 8678
rect 10039 8676 10063 8678
rect 10119 8676 10143 8678
rect 10199 8676 10205 8678
rect 9897 8667 10205 8676
rect 8852 8424 8904 8430
rect 9680 8424 9732 8430
rect 8904 8372 8984 8378
rect 8852 8366 8984 8372
rect 9680 8366 9732 8372
rect 8392 8356 8444 8362
rect 8864 8350 8984 8366
rect 8392 8298 8444 8304
rect 8404 6866 8432 8298
rect 8540 8188 8848 8197
rect 8540 8186 8546 8188
rect 8602 8186 8626 8188
rect 8682 8186 8706 8188
rect 8762 8186 8786 8188
rect 8842 8186 8848 8188
rect 8602 8134 8604 8186
rect 8784 8134 8786 8186
rect 8540 8132 8546 8134
rect 8602 8132 8626 8134
rect 8682 8132 8706 8134
rect 8762 8132 8786 8134
rect 8842 8132 8848 8134
rect 8540 8123 8848 8132
rect 8956 8090 8984 8350
rect 9036 8356 9088 8362
rect 9036 8298 9088 8304
rect 9496 8356 9548 8362
rect 9496 8298 9548 8304
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8944 7948 8996 7954
rect 8944 7890 8996 7896
rect 8956 7342 8984 7890
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 8540 7100 8848 7109
rect 8540 7098 8546 7100
rect 8602 7098 8626 7100
rect 8682 7098 8706 7100
rect 8762 7098 8786 7100
rect 8842 7098 8848 7100
rect 8602 7046 8604 7098
rect 8784 7046 8786 7098
rect 8540 7044 8546 7046
rect 8602 7044 8626 7046
rect 8682 7044 8706 7046
rect 8762 7044 8786 7046
rect 8842 7044 8848 7046
rect 8540 7035 8848 7044
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8392 6384 8444 6390
rect 8392 6326 8444 6332
rect 8850 6352 8906 6361
rect 8300 5840 8352 5846
rect 7838 5808 7894 5817
rect 7748 5772 7800 5778
rect 8300 5782 8352 5788
rect 8404 5778 8432 6326
rect 8850 6287 8906 6296
rect 8864 6254 8892 6287
rect 8852 6248 8904 6254
rect 8852 6190 8904 6196
rect 8540 6012 8848 6021
rect 8540 6010 8546 6012
rect 8602 6010 8626 6012
rect 8682 6010 8706 6012
rect 8762 6010 8786 6012
rect 8842 6010 8848 6012
rect 8602 5958 8604 6010
rect 8784 5958 8786 6010
rect 8540 5956 8546 5958
rect 8602 5956 8626 5958
rect 8682 5956 8706 5958
rect 8762 5956 8786 5958
rect 8842 5956 8848 5958
rect 8540 5947 8848 5956
rect 8956 5778 8984 7278
rect 9048 6458 9076 8298
rect 9312 8288 9364 8294
rect 9312 8230 9364 8236
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9140 7002 9168 7822
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 9232 7410 9260 7686
rect 9324 7546 9352 8230
rect 9404 7948 9456 7954
rect 9404 7890 9456 7896
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 9140 5914 9168 6190
rect 9232 5914 9260 7142
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 7838 5743 7894 5752
rect 8392 5772 8444 5778
rect 7748 5714 7800 5720
rect 8392 5714 8444 5720
rect 8944 5772 8996 5778
rect 8944 5714 8996 5720
rect 9416 5642 9444 7890
rect 9508 6322 9536 8298
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9600 6866 9628 7686
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9692 6662 9720 8366
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 9784 7206 9812 7822
rect 9897 7644 10205 7653
rect 9897 7642 9903 7644
rect 9959 7642 9983 7644
rect 10039 7642 10063 7644
rect 10119 7642 10143 7644
rect 10199 7642 10205 7644
rect 9959 7590 9961 7642
rect 10141 7590 10143 7642
rect 9897 7588 9903 7590
rect 9959 7588 9983 7590
rect 10039 7588 10063 7590
rect 10119 7588 10143 7590
rect 10199 7588 10205 7590
rect 9897 7579 10205 7588
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9692 6254 9720 6598
rect 9897 6556 10205 6565
rect 9897 6554 9903 6556
rect 9959 6554 9983 6556
rect 10039 6554 10063 6556
rect 10119 6554 10143 6556
rect 10199 6554 10205 6556
rect 9959 6502 9961 6554
rect 10141 6502 10143 6554
rect 9897 6500 9903 6502
rect 9959 6500 9983 6502
rect 10039 6500 10063 6502
rect 10119 6500 10143 6502
rect 10199 6500 10205 6502
rect 9897 6491 10205 6500
rect 10244 6458 10272 8910
rect 10336 8430 10364 9046
rect 10428 9042 10456 9318
rect 10416 9036 10468 9042
rect 10416 8978 10468 8984
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 10324 8424 10376 8430
rect 10324 8366 10376 8372
rect 10428 8022 10456 8774
rect 10520 8090 10548 9998
rect 10600 9648 10652 9654
rect 10600 9590 10652 9596
rect 10612 8090 10640 9590
rect 11072 9110 11100 10542
rect 11060 9104 11112 9110
rect 11060 9046 11112 9052
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10416 8016 10468 8022
rect 10416 7958 10468 7964
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 9680 6248 9732 6254
rect 9680 6190 9732 6196
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9508 5778 9536 6054
rect 9876 5778 9904 6394
rect 10324 6180 10376 6186
rect 10324 6122 10376 6128
rect 10232 5840 10284 5846
rect 10232 5782 10284 5788
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9864 5772 9916 5778
rect 9864 5714 9916 5720
rect 9404 5636 9456 5642
rect 9404 5578 9456 5584
rect 1755 5468 2063 5477
rect 1755 5466 1761 5468
rect 1817 5466 1841 5468
rect 1897 5466 1921 5468
rect 1977 5466 2001 5468
rect 2057 5466 2063 5468
rect 1817 5414 1819 5466
rect 1999 5414 2001 5466
rect 1755 5412 1761 5414
rect 1817 5412 1841 5414
rect 1897 5412 1921 5414
rect 1977 5412 2001 5414
rect 2057 5412 2063 5414
rect 1755 5403 2063 5412
rect 4469 5468 4777 5477
rect 4469 5466 4475 5468
rect 4531 5466 4555 5468
rect 4611 5466 4635 5468
rect 4691 5466 4715 5468
rect 4771 5466 4777 5468
rect 4531 5414 4533 5466
rect 4713 5414 4715 5466
rect 4469 5412 4475 5414
rect 4531 5412 4555 5414
rect 4611 5412 4635 5414
rect 4691 5412 4715 5414
rect 4771 5412 4777 5414
rect 4469 5403 4777 5412
rect 7183 5468 7491 5477
rect 7183 5466 7189 5468
rect 7245 5466 7269 5468
rect 7325 5466 7349 5468
rect 7405 5466 7429 5468
rect 7485 5466 7491 5468
rect 7245 5414 7247 5466
rect 7427 5414 7429 5466
rect 7183 5412 7189 5414
rect 7245 5412 7269 5414
rect 7325 5412 7349 5414
rect 7405 5412 7429 5414
rect 7485 5412 7491 5414
rect 7183 5403 7491 5412
rect 3112 4924 3420 4933
rect 3112 4922 3118 4924
rect 3174 4922 3198 4924
rect 3254 4922 3278 4924
rect 3334 4922 3358 4924
rect 3414 4922 3420 4924
rect 3174 4870 3176 4922
rect 3356 4870 3358 4922
rect 3112 4868 3118 4870
rect 3174 4868 3198 4870
rect 3254 4868 3278 4870
rect 3334 4868 3358 4870
rect 3414 4868 3420 4870
rect 3112 4859 3420 4868
rect 5826 4924 6134 4933
rect 5826 4922 5832 4924
rect 5888 4922 5912 4924
rect 5968 4922 5992 4924
rect 6048 4922 6072 4924
rect 6128 4922 6134 4924
rect 5888 4870 5890 4922
rect 6070 4870 6072 4922
rect 5826 4868 5832 4870
rect 5888 4868 5912 4870
rect 5968 4868 5992 4870
rect 6048 4868 6072 4870
rect 6128 4868 6134 4870
rect 5826 4859 6134 4868
rect 8540 4924 8848 4933
rect 8540 4922 8546 4924
rect 8602 4922 8626 4924
rect 8682 4922 8706 4924
rect 8762 4922 8786 4924
rect 8842 4922 8848 4924
rect 8602 4870 8604 4922
rect 8784 4870 8786 4922
rect 8540 4868 8546 4870
rect 8602 4868 8626 4870
rect 8682 4868 8706 4870
rect 8762 4868 8786 4870
rect 8842 4868 8848 4870
rect 8540 4859 8848 4868
rect 9508 4690 9536 5714
rect 9897 5468 10205 5477
rect 9897 5466 9903 5468
rect 9959 5466 9983 5468
rect 10039 5466 10063 5468
rect 10119 5466 10143 5468
rect 10199 5466 10205 5468
rect 9959 5414 9961 5466
rect 10141 5414 10143 5466
rect 9897 5412 9903 5414
rect 9959 5412 9983 5414
rect 10039 5412 10063 5414
rect 10119 5412 10143 5414
rect 10199 5412 10205 5414
rect 9897 5403 10205 5412
rect 10244 5302 10272 5782
rect 10336 5370 10364 6122
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10232 5296 10284 5302
rect 10232 5238 10284 5244
rect 10336 4758 10364 5306
rect 10428 5166 10456 7958
rect 10796 7410 10824 8910
rect 10968 8424 11020 8430
rect 10968 8366 11020 8372
rect 10980 8294 11008 8366
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 10980 7818 11008 8230
rect 11164 7886 11192 11342
rect 11254 10364 11562 10373
rect 11254 10362 11260 10364
rect 11316 10362 11340 10364
rect 11396 10362 11420 10364
rect 11476 10362 11500 10364
rect 11556 10362 11562 10364
rect 11316 10310 11318 10362
rect 11498 10310 11500 10362
rect 11254 10308 11260 10310
rect 11316 10308 11340 10310
rect 11396 10308 11420 10310
rect 11476 10308 11500 10310
rect 11556 10308 11562 10310
rect 11254 10299 11562 10308
rect 11254 9276 11562 9285
rect 11254 9274 11260 9276
rect 11316 9274 11340 9276
rect 11396 9274 11420 9276
rect 11476 9274 11500 9276
rect 11556 9274 11562 9276
rect 11316 9222 11318 9274
rect 11498 9222 11500 9274
rect 11254 9220 11260 9222
rect 11316 9220 11340 9222
rect 11396 9220 11420 9222
rect 11476 9220 11500 9222
rect 11556 9220 11562 9222
rect 11254 9211 11562 9220
rect 11254 8188 11562 8197
rect 11254 8186 11260 8188
rect 11316 8186 11340 8188
rect 11396 8186 11420 8188
rect 11476 8186 11500 8188
rect 11556 8186 11562 8188
rect 11316 8134 11318 8186
rect 11498 8134 11500 8186
rect 11254 8132 11260 8134
rect 11316 8132 11340 8134
rect 11396 8132 11420 8134
rect 11476 8132 11500 8134
rect 11556 8132 11562 8134
rect 11254 8123 11562 8132
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 10968 7812 11020 7818
rect 10968 7754 11020 7760
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 10520 5642 10548 7278
rect 10692 7200 10744 7206
rect 10692 7142 10744 7148
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10508 5636 10560 5642
rect 10508 5578 10560 5584
rect 10612 5370 10640 5646
rect 10600 5364 10652 5370
rect 10600 5306 10652 5312
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 10324 4752 10376 4758
rect 10324 4694 10376 4700
rect 10704 4690 10732 7142
rect 10796 7002 10824 7346
rect 10784 6996 10836 7002
rect 10784 6938 10836 6944
rect 10796 6338 10824 6938
rect 10796 6310 10916 6338
rect 10784 6180 10836 6186
rect 10784 6122 10836 6128
rect 10796 4826 10824 6122
rect 10888 5914 10916 6310
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10980 5098 11008 7754
rect 11254 7100 11562 7109
rect 11254 7098 11260 7100
rect 11316 7098 11340 7100
rect 11396 7098 11420 7100
rect 11476 7098 11500 7100
rect 11556 7098 11562 7100
rect 11316 7046 11318 7098
rect 11498 7046 11500 7098
rect 11254 7044 11260 7046
rect 11316 7044 11340 7046
rect 11396 7044 11420 7046
rect 11476 7044 11500 7046
rect 11556 7044 11562 7046
rect 11254 7035 11562 7044
rect 11254 6012 11562 6021
rect 11254 6010 11260 6012
rect 11316 6010 11340 6012
rect 11396 6010 11420 6012
rect 11476 6010 11500 6012
rect 11556 6010 11562 6012
rect 11316 5958 11318 6010
rect 11498 5958 11500 6010
rect 11254 5956 11260 5958
rect 11316 5956 11340 5958
rect 11396 5956 11420 5958
rect 11476 5956 11500 5958
rect 11556 5956 11562 5958
rect 11254 5947 11562 5956
rect 10968 5092 11020 5098
rect 10968 5034 11020 5040
rect 11254 4924 11562 4933
rect 11254 4922 11260 4924
rect 11316 4922 11340 4924
rect 11396 4922 11420 4924
rect 11476 4922 11500 4924
rect 11556 4922 11562 4924
rect 11316 4870 11318 4922
rect 11498 4870 11500 4922
rect 11254 4868 11260 4870
rect 11316 4868 11340 4870
rect 11396 4868 11420 4870
rect 11476 4868 11500 4870
rect 11556 4868 11562 4870
rect 11254 4859 11562 4868
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 10692 4684 10744 4690
rect 10692 4626 10744 4632
rect 1755 4380 2063 4389
rect 1755 4378 1761 4380
rect 1817 4378 1841 4380
rect 1897 4378 1921 4380
rect 1977 4378 2001 4380
rect 2057 4378 2063 4380
rect 1817 4326 1819 4378
rect 1999 4326 2001 4378
rect 1755 4324 1761 4326
rect 1817 4324 1841 4326
rect 1897 4324 1921 4326
rect 1977 4324 2001 4326
rect 2057 4324 2063 4326
rect 1755 4315 2063 4324
rect 4469 4380 4777 4389
rect 4469 4378 4475 4380
rect 4531 4378 4555 4380
rect 4611 4378 4635 4380
rect 4691 4378 4715 4380
rect 4771 4378 4777 4380
rect 4531 4326 4533 4378
rect 4713 4326 4715 4378
rect 4469 4324 4475 4326
rect 4531 4324 4555 4326
rect 4611 4324 4635 4326
rect 4691 4324 4715 4326
rect 4771 4324 4777 4326
rect 4469 4315 4777 4324
rect 7183 4380 7491 4389
rect 7183 4378 7189 4380
rect 7245 4378 7269 4380
rect 7325 4378 7349 4380
rect 7405 4378 7429 4380
rect 7485 4378 7491 4380
rect 7245 4326 7247 4378
rect 7427 4326 7429 4378
rect 7183 4324 7189 4326
rect 7245 4324 7269 4326
rect 7325 4324 7349 4326
rect 7405 4324 7429 4326
rect 7485 4324 7491 4326
rect 7183 4315 7491 4324
rect 9897 4380 10205 4389
rect 9897 4378 9903 4380
rect 9959 4378 9983 4380
rect 10039 4378 10063 4380
rect 10119 4378 10143 4380
rect 10199 4378 10205 4380
rect 9959 4326 9961 4378
rect 10141 4326 10143 4378
rect 9897 4324 9903 4326
rect 9959 4324 9983 4326
rect 10039 4324 10063 4326
rect 10119 4324 10143 4326
rect 10199 4324 10205 4326
rect 9897 4315 10205 4324
rect 3112 3836 3420 3845
rect 3112 3834 3118 3836
rect 3174 3834 3198 3836
rect 3254 3834 3278 3836
rect 3334 3834 3358 3836
rect 3414 3834 3420 3836
rect 3174 3782 3176 3834
rect 3356 3782 3358 3834
rect 3112 3780 3118 3782
rect 3174 3780 3198 3782
rect 3254 3780 3278 3782
rect 3334 3780 3358 3782
rect 3414 3780 3420 3782
rect 3112 3771 3420 3780
rect 5826 3836 6134 3845
rect 5826 3834 5832 3836
rect 5888 3834 5912 3836
rect 5968 3834 5992 3836
rect 6048 3834 6072 3836
rect 6128 3834 6134 3836
rect 5888 3782 5890 3834
rect 6070 3782 6072 3834
rect 5826 3780 5832 3782
rect 5888 3780 5912 3782
rect 5968 3780 5992 3782
rect 6048 3780 6072 3782
rect 6128 3780 6134 3782
rect 5826 3771 6134 3780
rect 8540 3836 8848 3845
rect 8540 3834 8546 3836
rect 8602 3834 8626 3836
rect 8682 3834 8706 3836
rect 8762 3834 8786 3836
rect 8842 3834 8848 3836
rect 8602 3782 8604 3834
rect 8784 3782 8786 3834
rect 8540 3780 8546 3782
rect 8602 3780 8626 3782
rect 8682 3780 8706 3782
rect 8762 3780 8786 3782
rect 8842 3780 8848 3782
rect 8540 3771 8848 3780
rect 11254 3836 11562 3845
rect 11254 3834 11260 3836
rect 11316 3834 11340 3836
rect 11396 3834 11420 3836
rect 11476 3834 11500 3836
rect 11556 3834 11562 3836
rect 11316 3782 11318 3834
rect 11498 3782 11500 3834
rect 11254 3780 11260 3782
rect 11316 3780 11340 3782
rect 11396 3780 11420 3782
rect 11476 3780 11500 3782
rect 11556 3780 11562 3782
rect 11254 3771 11562 3780
rect 1755 3292 2063 3301
rect 1755 3290 1761 3292
rect 1817 3290 1841 3292
rect 1897 3290 1921 3292
rect 1977 3290 2001 3292
rect 2057 3290 2063 3292
rect 1817 3238 1819 3290
rect 1999 3238 2001 3290
rect 1755 3236 1761 3238
rect 1817 3236 1841 3238
rect 1897 3236 1921 3238
rect 1977 3236 2001 3238
rect 2057 3236 2063 3238
rect 1755 3227 2063 3236
rect 4469 3292 4777 3301
rect 4469 3290 4475 3292
rect 4531 3290 4555 3292
rect 4611 3290 4635 3292
rect 4691 3290 4715 3292
rect 4771 3290 4777 3292
rect 4531 3238 4533 3290
rect 4713 3238 4715 3290
rect 4469 3236 4475 3238
rect 4531 3236 4555 3238
rect 4611 3236 4635 3238
rect 4691 3236 4715 3238
rect 4771 3236 4777 3238
rect 4469 3227 4777 3236
rect 7183 3292 7491 3301
rect 7183 3290 7189 3292
rect 7245 3290 7269 3292
rect 7325 3290 7349 3292
rect 7405 3290 7429 3292
rect 7485 3290 7491 3292
rect 7245 3238 7247 3290
rect 7427 3238 7429 3290
rect 7183 3236 7189 3238
rect 7245 3236 7269 3238
rect 7325 3236 7349 3238
rect 7405 3236 7429 3238
rect 7485 3236 7491 3238
rect 7183 3227 7491 3236
rect 9897 3292 10205 3301
rect 9897 3290 9903 3292
rect 9959 3290 9983 3292
rect 10039 3290 10063 3292
rect 10119 3290 10143 3292
rect 10199 3290 10205 3292
rect 9959 3238 9961 3290
rect 10141 3238 10143 3290
rect 9897 3236 9903 3238
rect 9959 3236 9983 3238
rect 10039 3236 10063 3238
rect 10119 3236 10143 3238
rect 10199 3236 10205 3238
rect 9897 3227 10205 3236
rect 3112 2748 3420 2757
rect 3112 2746 3118 2748
rect 3174 2746 3198 2748
rect 3254 2746 3278 2748
rect 3334 2746 3358 2748
rect 3414 2746 3420 2748
rect 3174 2694 3176 2746
rect 3356 2694 3358 2746
rect 3112 2692 3118 2694
rect 3174 2692 3198 2694
rect 3254 2692 3278 2694
rect 3334 2692 3358 2694
rect 3414 2692 3420 2694
rect 3112 2683 3420 2692
rect 5826 2748 6134 2757
rect 5826 2746 5832 2748
rect 5888 2746 5912 2748
rect 5968 2746 5992 2748
rect 6048 2746 6072 2748
rect 6128 2746 6134 2748
rect 5888 2694 5890 2746
rect 6070 2694 6072 2746
rect 5826 2692 5832 2694
rect 5888 2692 5912 2694
rect 5968 2692 5992 2694
rect 6048 2692 6072 2694
rect 6128 2692 6134 2694
rect 5826 2683 6134 2692
rect 8540 2748 8848 2757
rect 8540 2746 8546 2748
rect 8602 2746 8626 2748
rect 8682 2746 8706 2748
rect 8762 2746 8786 2748
rect 8842 2746 8848 2748
rect 8602 2694 8604 2746
rect 8784 2694 8786 2746
rect 8540 2692 8546 2694
rect 8602 2692 8626 2694
rect 8682 2692 8706 2694
rect 8762 2692 8786 2694
rect 8842 2692 8848 2694
rect 8540 2683 8848 2692
rect 11254 2748 11562 2757
rect 11254 2746 11260 2748
rect 11316 2746 11340 2748
rect 11396 2746 11420 2748
rect 11476 2746 11500 2748
rect 11556 2746 11562 2748
rect 11316 2694 11318 2746
rect 11498 2694 11500 2746
rect 11254 2692 11260 2694
rect 11316 2692 11340 2694
rect 11396 2692 11420 2694
rect 11476 2692 11500 2694
rect 11556 2692 11562 2694
rect 11254 2683 11562 2692
rect 1755 2204 2063 2213
rect 1755 2202 1761 2204
rect 1817 2202 1841 2204
rect 1897 2202 1921 2204
rect 1977 2202 2001 2204
rect 2057 2202 2063 2204
rect 1817 2150 1819 2202
rect 1999 2150 2001 2202
rect 1755 2148 1761 2150
rect 1817 2148 1841 2150
rect 1897 2148 1921 2150
rect 1977 2148 2001 2150
rect 2057 2148 2063 2150
rect 1755 2139 2063 2148
rect 4469 2204 4777 2213
rect 4469 2202 4475 2204
rect 4531 2202 4555 2204
rect 4611 2202 4635 2204
rect 4691 2202 4715 2204
rect 4771 2202 4777 2204
rect 4531 2150 4533 2202
rect 4713 2150 4715 2202
rect 4469 2148 4475 2150
rect 4531 2148 4555 2150
rect 4611 2148 4635 2150
rect 4691 2148 4715 2150
rect 4771 2148 4777 2150
rect 4469 2139 4777 2148
rect 7183 2204 7491 2213
rect 7183 2202 7189 2204
rect 7245 2202 7269 2204
rect 7325 2202 7349 2204
rect 7405 2202 7429 2204
rect 7485 2202 7491 2204
rect 7245 2150 7247 2202
rect 7427 2150 7429 2202
rect 7183 2148 7189 2150
rect 7245 2148 7269 2150
rect 7325 2148 7349 2150
rect 7405 2148 7429 2150
rect 7485 2148 7491 2150
rect 7183 2139 7491 2148
rect 9897 2204 10205 2213
rect 9897 2202 9903 2204
rect 9959 2202 9983 2204
rect 10039 2202 10063 2204
rect 10119 2202 10143 2204
rect 10199 2202 10205 2204
rect 9959 2150 9961 2202
rect 10141 2150 10143 2202
rect 9897 2148 9903 2150
rect 9959 2148 9983 2150
rect 10039 2148 10063 2150
rect 10119 2148 10143 2150
rect 10199 2148 10205 2150
rect 9897 2139 10205 2148
rect 3112 1660 3420 1669
rect 3112 1658 3118 1660
rect 3174 1658 3198 1660
rect 3254 1658 3278 1660
rect 3334 1658 3358 1660
rect 3414 1658 3420 1660
rect 3174 1606 3176 1658
rect 3356 1606 3358 1658
rect 3112 1604 3118 1606
rect 3174 1604 3198 1606
rect 3254 1604 3278 1606
rect 3334 1604 3358 1606
rect 3414 1604 3420 1606
rect 3112 1595 3420 1604
rect 5826 1660 6134 1669
rect 5826 1658 5832 1660
rect 5888 1658 5912 1660
rect 5968 1658 5992 1660
rect 6048 1658 6072 1660
rect 6128 1658 6134 1660
rect 5888 1606 5890 1658
rect 6070 1606 6072 1658
rect 5826 1604 5832 1606
rect 5888 1604 5912 1606
rect 5968 1604 5992 1606
rect 6048 1604 6072 1606
rect 6128 1604 6134 1606
rect 5826 1595 6134 1604
rect 8540 1660 8848 1669
rect 8540 1658 8546 1660
rect 8602 1658 8626 1660
rect 8682 1658 8706 1660
rect 8762 1658 8786 1660
rect 8842 1658 8848 1660
rect 8602 1606 8604 1658
rect 8784 1606 8786 1658
rect 8540 1604 8546 1606
rect 8602 1604 8626 1606
rect 8682 1604 8706 1606
rect 8762 1604 8786 1606
rect 8842 1604 8848 1606
rect 8540 1595 8848 1604
rect 11254 1660 11562 1669
rect 11254 1658 11260 1660
rect 11316 1658 11340 1660
rect 11396 1658 11420 1660
rect 11476 1658 11500 1660
rect 11556 1658 11562 1660
rect 11316 1606 11318 1658
rect 11498 1606 11500 1658
rect 11254 1604 11260 1606
rect 11316 1604 11340 1606
rect 11396 1604 11420 1606
rect 11476 1604 11500 1606
rect 11556 1604 11562 1606
rect 11254 1595 11562 1604
rect 1755 1116 2063 1125
rect 1755 1114 1761 1116
rect 1817 1114 1841 1116
rect 1897 1114 1921 1116
rect 1977 1114 2001 1116
rect 2057 1114 2063 1116
rect 1817 1062 1819 1114
rect 1999 1062 2001 1114
rect 1755 1060 1761 1062
rect 1817 1060 1841 1062
rect 1897 1060 1921 1062
rect 1977 1060 2001 1062
rect 2057 1060 2063 1062
rect 1755 1051 2063 1060
rect 4469 1116 4777 1125
rect 4469 1114 4475 1116
rect 4531 1114 4555 1116
rect 4611 1114 4635 1116
rect 4691 1114 4715 1116
rect 4771 1114 4777 1116
rect 4531 1062 4533 1114
rect 4713 1062 4715 1114
rect 4469 1060 4475 1062
rect 4531 1060 4555 1062
rect 4611 1060 4635 1062
rect 4691 1060 4715 1062
rect 4771 1060 4777 1062
rect 4469 1051 4777 1060
rect 7183 1116 7491 1125
rect 7183 1114 7189 1116
rect 7245 1114 7269 1116
rect 7325 1114 7349 1116
rect 7405 1114 7429 1116
rect 7485 1114 7491 1116
rect 7245 1062 7247 1114
rect 7427 1062 7429 1114
rect 7183 1060 7189 1062
rect 7245 1060 7269 1062
rect 7325 1060 7349 1062
rect 7405 1060 7429 1062
rect 7485 1060 7491 1062
rect 7183 1051 7491 1060
rect 9897 1116 10205 1125
rect 9897 1114 9903 1116
rect 9959 1114 9983 1116
rect 10039 1114 10063 1116
rect 10119 1114 10143 1116
rect 10199 1114 10205 1116
rect 9959 1062 9961 1114
rect 10141 1062 10143 1114
rect 9897 1060 9903 1062
rect 9959 1060 9983 1062
rect 10039 1060 10063 1062
rect 10119 1060 10143 1062
rect 10199 1060 10205 1062
rect 9897 1051 10205 1060
rect 3112 572 3420 581
rect 3112 570 3118 572
rect 3174 570 3198 572
rect 3254 570 3278 572
rect 3334 570 3358 572
rect 3414 570 3420 572
rect 3174 518 3176 570
rect 3356 518 3358 570
rect 3112 516 3118 518
rect 3174 516 3198 518
rect 3254 516 3278 518
rect 3334 516 3358 518
rect 3414 516 3420 518
rect 3112 507 3420 516
rect 5826 572 6134 581
rect 5826 570 5832 572
rect 5888 570 5912 572
rect 5968 570 5992 572
rect 6048 570 6072 572
rect 6128 570 6134 572
rect 5888 518 5890 570
rect 6070 518 6072 570
rect 5826 516 5832 518
rect 5888 516 5912 518
rect 5968 516 5992 518
rect 6048 516 6072 518
rect 6128 516 6134 518
rect 5826 507 6134 516
rect 8540 572 8848 581
rect 8540 570 8546 572
rect 8602 570 8626 572
rect 8682 570 8706 572
rect 8762 570 8786 572
rect 8842 570 8848 572
rect 8602 518 8604 570
rect 8784 518 8786 570
rect 8540 516 8546 518
rect 8602 516 8626 518
rect 8682 516 8706 518
rect 8762 516 8786 518
rect 8842 516 8848 518
rect 8540 507 8848 516
rect 11254 572 11562 581
rect 11254 570 11260 572
rect 11316 570 11340 572
rect 11396 570 11420 572
rect 11476 570 11500 572
rect 11556 570 11562 572
rect 11316 518 11318 570
rect 11498 518 11500 570
rect 11254 516 11260 518
rect 11316 516 11340 518
rect 11396 516 11420 518
rect 11476 516 11500 518
rect 11556 516 11562 518
rect 11254 507 11562 516
<< via2 >>
rect 1761 10906 1817 10908
rect 1841 10906 1897 10908
rect 1921 10906 1977 10908
rect 2001 10906 2057 10908
rect 1761 10854 1807 10906
rect 1807 10854 1817 10906
rect 1841 10854 1871 10906
rect 1871 10854 1883 10906
rect 1883 10854 1897 10906
rect 1921 10854 1935 10906
rect 1935 10854 1947 10906
rect 1947 10854 1977 10906
rect 2001 10854 2011 10906
rect 2011 10854 2057 10906
rect 1761 10852 1817 10854
rect 1841 10852 1897 10854
rect 1921 10852 1977 10854
rect 2001 10852 2057 10854
rect 1214 9560 1270 9616
rect 1761 9818 1817 9820
rect 1841 9818 1897 9820
rect 1921 9818 1977 9820
rect 2001 9818 2057 9820
rect 1761 9766 1807 9818
rect 1807 9766 1817 9818
rect 1841 9766 1871 9818
rect 1871 9766 1883 9818
rect 1883 9766 1897 9818
rect 1921 9766 1935 9818
rect 1935 9766 1947 9818
rect 1947 9766 1977 9818
rect 2001 9766 2011 9818
rect 2011 9766 2057 9818
rect 1761 9764 1817 9766
rect 1841 9764 1897 9766
rect 1921 9764 1977 9766
rect 2001 9764 2057 9766
rect 3118 11450 3174 11452
rect 3198 11450 3254 11452
rect 3278 11450 3334 11452
rect 3358 11450 3414 11452
rect 3118 11398 3164 11450
rect 3164 11398 3174 11450
rect 3198 11398 3228 11450
rect 3228 11398 3240 11450
rect 3240 11398 3254 11450
rect 3278 11398 3292 11450
rect 3292 11398 3304 11450
rect 3304 11398 3334 11450
rect 3358 11398 3368 11450
rect 3368 11398 3414 11450
rect 3118 11396 3174 11398
rect 3198 11396 3254 11398
rect 3278 11396 3334 11398
rect 3358 11396 3414 11398
rect 5832 11450 5888 11452
rect 5912 11450 5968 11452
rect 5992 11450 6048 11452
rect 6072 11450 6128 11452
rect 5832 11398 5878 11450
rect 5878 11398 5888 11450
rect 5912 11398 5942 11450
rect 5942 11398 5954 11450
rect 5954 11398 5968 11450
rect 5992 11398 6006 11450
rect 6006 11398 6018 11450
rect 6018 11398 6048 11450
rect 6072 11398 6082 11450
rect 6082 11398 6128 11450
rect 5832 11396 5888 11398
rect 5912 11396 5968 11398
rect 5992 11396 6048 11398
rect 6072 11396 6128 11398
rect 1761 8730 1817 8732
rect 1841 8730 1897 8732
rect 1921 8730 1977 8732
rect 2001 8730 2057 8732
rect 1761 8678 1807 8730
rect 1807 8678 1817 8730
rect 1841 8678 1871 8730
rect 1871 8678 1883 8730
rect 1883 8678 1897 8730
rect 1921 8678 1935 8730
rect 1935 8678 1947 8730
rect 1947 8678 1977 8730
rect 2001 8678 2011 8730
rect 2011 8678 2057 8730
rect 1761 8676 1817 8678
rect 1841 8676 1897 8678
rect 1921 8676 1977 8678
rect 2001 8676 2057 8678
rect 4475 10906 4531 10908
rect 4555 10906 4611 10908
rect 4635 10906 4691 10908
rect 4715 10906 4771 10908
rect 4475 10854 4521 10906
rect 4521 10854 4531 10906
rect 4555 10854 4585 10906
rect 4585 10854 4597 10906
rect 4597 10854 4611 10906
rect 4635 10854 4649 10906
rect 4649 10854 4661 10906
rect 4661 10854 4691 10906
rect 4715 10854 4725 10906
rect 4725 10854 4771 10906
rect 4475 10852 4531 10854
rect 4555 10852 4611 10854
rect 4635 10852 4691 10854
rect 4715 10852 4771 10854
rect 3118 10362 3174 10364
rect 3198 10362 3254 10364
rect 3278 10362 3334 10364
rect 3358 10362 3414 10364
rect 3118 10310 3164 10362
rect 3164 10310 3174 10362
rect 3198 10310 3228 10362
rect 3228 10310 3240 10362
rect 3240 10310 3254 10362
rect 3278 10310 3292 10362
rect 3292 10310 3304 10362
rect 3304 10310 3334 10362
rect 3358 10310 3368 10362
rect 3368 10310 3414 10362
rect 3118 10308 3174 10310
rect 3198 10308 3254 10310
rect 3278 10308 3334 10310
rect 3358 10308 3414 10310
rect 3330 9560 3386 9616
rect 3054 9460 3056 9480
rect 3056 9460 3108 9480
rect 3108 9460 3110 9480
rect 3054 9424 3110 9460
rect 3118 9274 3174 9276
rect 3198 9274 3254 9276
rect 3278 9274 3334 9276
rect 3358 9274 3414 9276
rect 3118 9222 3164 9274
rect 3164 9222 3174 9274
rect 3198 9222 3228 9274
rect 3228 9222 3240 9274
rect 3240 9222 3254 9274
rect 3278 9222 3292 9274
rect 3292 9222 3304 9274
rect 3304 9222 3334 9274
rect 3358 9222 3368 9274
rect 3368 9222 3414 9274
rect 3118 9220 3174 9222
rect 3198 9220 3254 9222
rect 3278 9220 3334 9222
rect 3358 9220 3414 9222
rect 3118 8186 3174 8188
rect 3198 8186 3254 8188
rect 3278 8186 3334 8188
rect 3358 8186 3414 8188
rect 3118 8134 3164 8186
rect 3164 8134 3174 8186
rect 3198 8134 3228 8186
rect 3228 8134 3240 8186
rect 3240 8134 3254 8186
rect 3278 8134 3292 8186
rect 3292 8134 3304 8186
rect 3304 8134 3334 8186
rect 3358 8134 3368 8186
rect 3368 8134 3414 8186
rect 3118 8132 3174 8134
rect 3198 8132 3254 8134
rect 3278 8132 3334 8134
rect 3358 8132 3414 8134
rect 1761 7642 1817 7644
rect 1841 7642 1897 7644
rect 1921 7642 1977 7644
rect 2001 7642 2057 7644
rect 1761 7590 1807 7642
rect 1807 7590 1817 7642
rect 1841 7590 1871 7642
rect 1871 7590 1883 7642
rect 1883 7590 1897 7642
rect 1921 7590 1935 7642
rect 1935 7590 1947 7642
rect 1947 7590 1977 7642
rect 2001 7590 2011 7642
rect 2011 7590 2057 7642
rect 1761 7588 1817 7590
rect 1841 7588 1897 7590
rect 1921 7588 1977 7590
rect 2001 7588 2057 7590
rect 1761 6554 1817 6556
rect 1841 6554 1897 6556
rect 1921 6554 1977 6556
rect 2001 6554 2057 6556
rect 1761 6502 1807 6554
rect 1807 6502 1817 6554
rect 1841 6502 1871 6554
rect 1871 6502 1883 6554
rect 1883 6502 1897 6554
rect 1921 6502 1935 6554
rect 1935 6502 1947 6554
rect 1947 6502 1977 6554
rect 2001 6502 2011 6554
rect 2011 6502 2057 6554
rect 1761 6500 1817 6502
rect 1841 6500 1897 6502
rect 1921 6500 1977 6502
rect 2001 6500 2057 6502
rect 3118 7098 3174 7100
rect 3198 7098 3254 7100
rect 3278 7098 3334 7100
rect 3358 7098 3414 7100
rect 3118 7046 3164 7098
rect 3164 7046 3174 7098
rect 3198 7046 3228 7098
rect 3228 7046 3240 7098
rect 3240 7046 3254 7098
rect 3278 7046 3292 7098
rect 3292 7046 3304 7098
rect 3304 7046 3334 7098
rect 3358 7046 3368 7098
rect 3368 7046 3414 7098
rect 3118 7044 3174 7046
rect 3198 7044 3254 7046
rect 3278 7044 3334 7046
rect 3358 7044 3414 7046
rect 4475 9818 4531 9820
rect 4555 9818 4611 9820
rect 4635 9818 4691 9820
rect 4715 9818 4771 9820
rect 4475 9766 4521 9818
rect 4521 9766 4531 9818
rect 4555 9766 4585 9818
rect 4585 9766 4597 9818
rect 4597 9766 4611 9818
rect 4635 9766 4649 9818
rect 4649 9766 4661 9818
rect 4661 9766 4691 9818
rect 4715 9766 4725 9818
rect 4725 9766 4771 9818
rect 4475 9764 4531 9766
rect 4555 9764 4611 9766
rect 4635 9764 4691 9766
rect 4715 9764 4771 9766
rect 4475 8730 4531 8732
rect 4555 8730 4611 8732
rect 4635 8730 4691 8732
rect 4715 8730 4771 8732
rect 4475 8678 4521 8730
rect 4521 8678 4531 8730
rect 4555 8678 4585 8730
rect 4585 8678 4597 8730
rect 4597 8678 4611 8730
rect 4635 8678 4649 8730
rect 4649 8678 4661 8730
rect 4661 8678 4691 8730
rect 4715 8678 4725 8730
rect 4725 8678 4771 8730
rect 4475 8676 4531 8678
rect 4555 8676 4611 8678
rect 4635 8676 4691 8678
rect 4715 8676 4771 8678
rect 5446 9968 5502 10024
rect 5262 9444 5318 9480
rect 5262 9424 5264 9444
rect 5264 9424 5316 9444
rect 5316 9424 5318 9444
rect 5832 10362 5888 10364
rect 5912 10362 5968 10364
rect 5992 10362 6048 10364
rect 6072 10362 6128 10364
rect 5832 10310 5878 10362
rect 5878 10310 5888 10362
rect 5912 10310 5942 10362
rect 5942 10310 5954 10362
rect 5954 10310 5968 10362
rect 5992 10310 6006 10362
rect 6006 10310 6018 10362
rect 6018 10310 6048 10362
rect 6072 10310 6082 10362
rect 6082 10310 6128 10362
rect 5832 10308 5888 10310
rect 5912 10308 5968 10310
rect 5992 10308 6048 10310
rect 6072 10308 6128 10310
rect 7189 10906 7245 10908
rect 7269 10906 7325 10908
rect 7349 10906 7405 10908
rect 7429 10906 7485 10908
rect 7189 10854 7235 10906
rect 7235 10854 7245 10906
rect 7269 10854 7299 10906
rect 7299 10854 7311 10906
rect 7311 10854 7325 10906
rect 7349 10854 7363 10906
rect 7363 10854 7375 10906
rect 7375 10854 7405 10906
rect 7429 10854 7439 10906
rect 7439 10854 7485 10906
rect 7189 10852 7245 10854
rect 7269 10852 7325 10854
rect 7349 10852 7405 10854
rect 7429 10852 7485 10854
rect 8546 11450 8602 11452
rect 8626 11450 8682 11452
rect 8706 11450 8762 11452
rect 8786 11450 8842 11452
rect 8546 11398 8592 11450
rect 8592 11398 8602 11450
rect 8626 11398 8656 11450
rect 8656 11398 8668 11450
rect 8668 11398 8682 11450
rect 8706 11398 8720 11450
rect 8720 11398 8732 11450
rect 8732 11398 8762 11450
rect 8786 11398 8796 11450
rect 8796 11398 8842 11450
rect 8546 11396 8602 11398
rect 8626 11396 8682 11398
rect 8706 11396 8762 11398
rect 8786 11396 8842 11398
rect 7189 9818 7245 9820
rect 7269 9818 7325 9820
rect 7349 9818 7405 9820
rect 7429 9818 7485 9820
rect 7189 9766 7235 9818
rect 7235 9766 7245 9818
rect 7269 9766 7299 9818
rect 7299 9766 7311 9818
rect 7311 9766 7325 9818
rect 7349 9766 7363 9818
rect 7363 9766 7375 9818
rect 7375 9766 7405 9818
rect 7429 9766 7439 9818
rect 7439 9766 7485 9818
rect 7189 9764 7245 9766
rect 7269 9764 7325 9766
rect 7349 9764 7405 9766
rect 7429 9764 7485 9766
rect 6826 9424 6882 9480
rect 7286 9424 7342 9480
rect 5832 9274 5888 9276
rect 5912 9274 5968 9276
rect 5992 9274 6048 9276
rect 6072 9274 6128 9276
rect 5832 9222 5878 9274
rect 5878 9222 5888 9274
rect 5912 9222 5942 9274
rect 5942 9222 5954 9274
rect 5954 9222 5968 9274
rect 5992 9222 6006 9274
rect 6006 9222 6018 9274
rect 6018 9222 6048 9274
rect 6072 9222 6082 9274
rect 6082 9222 6128 9274
rect 5832 9220 5888 9222
rect 5912 9220 5968 9222
rect 5992 9220 6048 9222
rect 6072 9220 6128 9222
rect 4475 7642 4531 7644
rect 4555 7642 4611 7644
rect 4635 7642 4691 7644
rect 4715 7642 4771 7644
rect 4475 7590 4521 7642
rect 4521 7590 4531 7642
rect 4555 7590 4585 7642
rect 4585 7590 4597 7642
rect 4597 7590 4611 7642
rect 4635 7590 4649 7642
rect 4649 7590 4661 7642
rect 4661 7590 4691 7642
rect 4715 7590 4725 7642
rect 4725 7590 4771 7642
rect 4475 7588 4531 7590
rect 4555 7588 4611 7590
rect 4635 7588 4691 7590
rect 4715 7588 4771 7590
rect 4475 6554 4531 6556
rect 4555 6554 4611 6556
rect 4635 6554 4691 6556
rect 4715 6554 4771 6556
rect 4475 6502 4521 6554
rect 4521 6502 4531 6554
rect 4555 6502 4585 6554
rect 4585 6502 4597 6554
rect 4597 6502 4611 6554
rect 4635 6502 4649 6554
rect 4649 6502 4661 6554
rect 4661 6502 4691 6554
rect 4715 6502 4725 6554
rect 4725 6502 4771 6554
rect 4475 6500 4531 6502
rect 4555 6500 4611 6502
rect 4635 6500 4691 6502
rect 4715 6500 4771 6502
rect 5832 8186 5888 8188
rect 5912 8186 5968 8188
rect 5992 8186 6048 8188
rect 6072 8186 6128 8188
rect 5832 8134 5878 8186
rect 5878 8134 5888 8186
rect 5912 8134 5942 8186
rect 5942 8134 5954 8186
rect 5954 8134 5968 8186
rect 5992 8134 6006 8186
rect 6006 8134 6018 8186
rect 6018 8134 6048 8186
rect 6072 8134 6082 8186
rect 6082 8134 6128 8186
rect 5832 8132 5888 8134
rect 5912 8132 5968 8134
rect 5992 8132 6048 8134
rect 6072 8132 6128 8134
rect 5832 7098 5888 7100
rect 5912 7098 5968 7100
rect 5992 7098 6048 7100
rect 6072 7098 6128 7100
rect 5832 7046 5878 7098
rect 5878 7046 5888 7098
rect 5912 7046 5942 7098
rect 5942 7046 5954 7098
rect 5954 7046 5968 7098
rect 5992 7046 6006 7098
rect 6006 7046 6018 7098
rect 6018 7046 6048 7098
rect 6072 7046 6082 7098
rect 6082 7046 6128 7098
rect 5832 7044 5888 7046
rect 5912 7044 5968 7046
rect 5992 7044 6048 7046
rect 6072 7044 6128 7046
rect 7189 8730 7245 8732
rect 7269 8730 7325 8732
rect 7349 8730 7405 8732
rect 7429 8730 7485 8732
rect 7189 8678 7235 8730
rect 7235 8678 7245 8730
rect 7269 8678 7299 8730
rect 7299 8678 7311 8730
rect 7311 8678 7325 8730
rect 7349 8678 7363 8730
rect 7363 8678 7375 8730
rect 7375 8678 7405 8730
rect 7429 8678 7439 8730
rect 7439 8678 7485 8730
rect 7189 8676 7245 8678
rect 7269 8676 7325 8678
rect 7349 8676 7405 8678
rect 7429 8676 7485 8678
rect 7189 7642 7245 7644
rect 7269 7642 7325 7644
rect 7349 7642 7405 7644
rect 7429 7642 7485 7644
rect 7189 7590 7235 7642
rect 7235 7590 7245 7642
rect 7269 7590 7299 7642
rect 7299 7590 7311 7642
rect 7311 7590 7325 7642
rect 7349 7590 7363 7642
rect 7363 7590 7375 7642
rect 7375 7590 7405 7642
rect 7429 7590 7439 7642
rect 7439 7590 7485 7642
rect 7189 7588 7245 7590
rect 7269 7588 7325 7590
rect 7349 7588 7405 7590
rect 7429 7588 7485 7590
rect 7189 6554 7245 6556
rect 7269 6554 7325 6556
rect 7349 6554 7405 6556
rect 7429 6554 7485 6556
rect 7189 6502 7235 6554
rect 7235 6502 7245 6554
rect 7269 6502 7299 6554
rect 7299 6502 7311 6554
rect 7311 6502 7325 6554
rect 7349 6502 7363 6554
rect 7363 6502 7375 6554
rect 7375 6502 7405 6554
rect 7429 6502 7439 6554
rect 7439 6502 7485 6554
rect 7189 6500 7245 6502
rect 7269 6500 7325 6502
rect 7349 6500 7405 6502
rect 7429 6500 7485 6502
rect 3118 6010 3174 6012
rect 3198 6010 3254 6012
rect 3278 6010 3334 6012
rect 3358 6010 3414 6012
rect 3118 5958 3164 6010
rect 3164 5958 3174 6010
rect 3198 5958 3228 6010
rect 3228 5958 3240 6010
rect 3240 5958 3254 6010
rect 3278 5958 3292 6010
rect 3292 5958 3304 6010
rect 3304 5958 3334 6010
rect 3358 5958 3368 6010
rect 3368 5958 3414 6010
rect 3118 5956 3174 5958
rect 3198 5956 3254 5958
rect 3278 5956 3334 5958
rect 3358 5956 3414 5958
rect 5832 6010 5888 6012
rect 5912 6010 5968 6012
rect 5992 6010 6048 6012
rect 6072 6010 6128 6012
rect 5832 5958 5878 6010
rect 5878 5958 5888 6010
rect 5912 5958 5942 6010
rect 5942 5958 5954 6010
rect 5954 5958 5968 6010
rect 5992 5958 6006 6010
rect 6006 5958 6018 6010
rect 6018 5958 6048 6010
rect 6072 5958 6082 6010
rect 6082 5958 6128 6010
rect 5832 5956 5888 5958
rect 5912 5956 5968 5958
rect 5992 5956 6048 5958
rect 6072 5956 6128 5958
rect 8546 10362 8602 10364
rect 8626 10362 8682 10364
rect 8706 10362 8762 10364
rect 8786 10362 8842 10364
rect 8546 10310 8592 10362
rect 8592 10310 8602 10362
rect 8626 10310 8656 10362
rect 8656 10310 8668 10362
rect 8668 10310 8682 10362
rect 8706 10310 8720 10362
rect 8720 10310 8732 10362
rect 8732 10310 8762 10362
rect 8786 10310 8796 10362
rect 8796 10310 8842 10362
rect 8546 10308 8602 10310
rect 8626 10308 8682 10310
rect 8706 10308 8762 10310
rect 8786 10308 8842 10310
rect 9310 9560 9366 9616
rect 11260 11450 11316 11452
rect 11340 11450 11396 11452
rect 11420 11450 11476 11452
rect 11500 11450 11556 11452
rect 11260 11398 11306 11450
rect 11306 11398 11316 11450
rect 11340 11398 11370 11450
rect 11370 11398 11382 11450
rect 11382 11398 11396 11450
rect 11420 11398 11434 11450
rect 11434 11398 11446 11450
rect 11446 11398 11476 11450
rect 11500 11398 11510 11450
rect 11510 11398 11556 11450
rect 11260 11396 11316 11398
rect 11340 11396 11396 11398
rect 11420 11396 11476 11398
rect 11500 11396 11556 11398
rect 9903 10906 9959 10908
rect 9983 10906 10039 10908
rect 10063 10906 10119 10908
rect 10143 10906 10199 10908
rect 9903 10854 9949 10906
rect 9949 10854 9959 10906
rect 9983 10854 10013 10906
rect 10013 10854 10025 10906
rect 10025 10854 10039 10906
rect 10063 10854 10077 10906
rect 10077 10854 10089 10906
rect 10089 10854 10119 10906
rect 10143 10854 10153 10906
rect 10153 10854 10199 10906
rect 9903 10852 9959 10854
rect 9983 10852 10039 10854
rect 10063 10852 10119 10854
rect 10143 10852 10199 10854
rect 9770 9968 9826 10024
rect 8666 9460 8668 9480
rect 8668 9460 8720 9480
rect 8720 9460 8722 9480
rect 8666 9424 8722 9460
rect 8546 9274 8602 9276
rect 8626 9274 8682 9276
rect 8706 9274 8762 9276
rect 8786 9274 8842 9276
rect 8546 9222 8592 9274
rect 8592 9222 8602 9274
rect 8626 9222 8656 9274
rect 8656 9222 8668 9274
rect 8668 9222 8682 9274
rect 8706 9222 8720 9274
rect 8720 9222 8732 9274
rect 8732 9222 8762 9274
rect 8786 9222 8796 9274
rect 8796 9222 8842 9274
rect 8546 9220 8602 9222
rect 8626 9220 8682 9222
rect 8706 9220 8762 9222
rect 8786 9220 8842 9222
rect 9903 9818 9959 9820
rect 9983 9818 10039 9820
rect 10063 9818 10119 9820
rect 10143 9818 10199 9820
rect 9903 9766 9949 9818
rect 9949 9766 9959 9818
rect 9983 9766 10013 9818
rect 10013 9766 10025 9818
rect 10025 9766 10039 9818
rect 10063 9766 10077 9818
rect 10077 9766 10089 9818
rect 10089 9766 10119 9818
rect 10143 9766 10153 9818
rect 10153 9766 10199 9818
rect 9903 9764 9959 9766
rect 9983 9764 10039 9766
rect 10063 9764 10119 9766
rect 10143 9764 10199 9766
rect 9903 8730 9959 8732
rect 9983 8730 10039 8732
rect 10063 8730 10119 8732
rect 10143 8730 10199 8732
rect 9903 8678 9949 8730
rect 9949 8678 9959 8730
rect 9983 8678 10013 8730
rect 10013 8678 10025 8730
rect 10025 8678 10039 8730
rect 10063 8678 10077 8730
rect 10077 8678 10089 8730
rect 10089 8678 10119 8730
rect 10143 8678 10153 8730
rect 10153 8678 10199 8730
rect 9903 8676 9959 8678
rect 9983 8676 10039 8678
rect 10063 8676 10119 8678
rect 10143 8676 10199 8678
rect 8546 8186 8602 8188
rect 8626 8186 8682 8188
rect 8706 8186 8762 8188
rect 8786 8186 8842 8188
rect 8546 8134 8592 8186
rect 8592 8134 8602 8186
rect 8626 8134 8656 8186
rect 8656 8134 8668 8186
rect 8668 8134 8682 8186
rect 8706 8134 8720 8186
rect 8720 8134 8732 8186
rect 8732 8134 8762 8186
rect 8786 8134 8796 8186
rect 8796 8134 8842 8186
rect 8546 8132 8602 8134
rect 8626 8132 8682 8134
rect 8706 8132 8762 8134
rect 8786 8132 8842 8134
rect 8546 7098 8602 7100
rect 8626 7098 8682 7100
rect 8706 7098 8762 7100
rect 8786 7098 8842 7100
rect 8546 7046 8592 7098
rect 8592 7046 8602 7098
rect 8626 7046 8656 7098
rect 8656 7046 8668 7098
rect 8668 7046 8682 7098
rect 8706 7046 8720 7098
rect 8720 7046 8732 7098
rect 8732 7046 8762 7098
rect 8786 7046 8796 7098
rect 8796 7046 8842 7098
rect 8546 7044 8602 7046
rect 8626 7044 8682 7046
rect 8706 7044 8762 7046
rect 8786 7044 8842 7046
rect 7838 5752 7894 5808
rect 8850 6296 8906 6352
rect 8546 6010 8602 6012
rect 8626 6010 8682 6012
rect 8706 6010 8762 6012
rect 8786 6010 8842 6012
rect 8546 5958 8592 6010
rect 8592 5958 8602 6010
rect 8626 5958 8656 6010
rect 8656 5958 8668 6010
rect 8668 5958 8682 6010
rect 8706 5958 8720 6010
rect 8720 5958 8732 6010
rect 8732 5958 8762 6010
rect 8786 5958 8796 6010
rect 8796 5958 8842 6010
rect 8546 5956 8602 5958
rect 8626 5956 8682 5958
rect 8706 5956 8762 5958
rect 8786 5956 8842 5958
rect 9903 7642 9959 7644
rect 9983 7642 10039 7644
rect 10063 7642 10119 7644
rect 10143 7642 10199 7644
rect 9903 7590 9949 7642
rect 9949 7590 9959 7642
rect 9983 7590 10013 7642
rect 10013 7590 10025 7642
rect 10025 7590 10039 7642
rect 10063 7590 10077 7642
rect 10077 7590 10089 7642
rect 10089 7590 10119 7642
rect 10143 7590 10153 7642
rect 10153 7590 10199 7642
rect 9903 7588 9959 7590
rect 9983 7588 10039 7590
rect 10063 7588 10119 7590
rect 10143 7588 10199 7590
rect 9903 6554 9959 6556
rect 9983 6554 10039 6556
rect 10063 6554 10119 6556
rect 10143 6554 10199 6556
rect 9903 6502 9949 6554
rect 9949 6502 9959 6554
rect 9983 6502 10013 6554
rect 10013 6502 10025 6554
rect 10025 6502 10039 6554
rect 10063 6502 10077 6554
rect 10077 6502 10089 6554
rect 10089 6502 10119 6554
rect 10143 6502 10153 6554
rect 10153 6502 10199 6554
rect 9903 6500 9959 6502
rect 9983 6500 10039 6502
rect 10063 6500 10119 6502
rect 10143 6500 10199 6502
rect 1761 5466 1817 5468
rect 1841 5466 1897 5468
rect 1921 5466 1977 5468
rect 2001 5466 2057 5468
rect 1761 5414 1807 5466
rect 1807 5414 1817 5466
rect 1841 5414 1871 5466
rect 1871 5414 1883 5466
rect 1883 5414 1897 5466
rect 1921 5414 1935 5466
rect 1935 5414 1947 5466
rect 1947 5414 1977 5466
rect 2001 5414 2011 5466
rect 2011 5414 2057 5466
rect 1761 5412 1817 5414
rect 1841 5412 1897 5414
rect 1921 5412 1977 5414
rect 2001 5412 2057 5414
rect 4475 5466 4531 5468
rect 4555 5466 4611 5468
rect 4635 5466 4691 5468
rect 4715 5466 4771 5468
rect 4475 5414 4521 5466
rect 4521 5414 4531 5466
rect 4555 5414 4585 5466
rect 4585 5414 4597 5466
rect 4597 5414 4611 5466
rect 4635 5414 4649 5466
rect 4649 5414 4661 5466
rect 4661 5414 4691 5466
rect 4715 5414 4725 5466
rect 4725 5414 4771 5466
rect 4475 5412 4531 5414
rect 4555 5412 4611 5414
rect 4635 5412 4691 5414
rect 4715 5412 4771 5414
rect 7189 5466 7245 5468
rect 7269 5466 7325 5468
rect 7349 5466 7405 5468
rect 7429 5466 7485 5468
rect 7189 5414 7235 5466
rect 7235 5414 7245 5466
rect 7269 5414 7299 5466
rect 7299 5414 7311 5466
rect 7311 5414 7325 5466
rect 7349 5414 7363 5466
rect 7363 5414 7375 5466
rect 7375 5414 7405 5466
rect 7429 5414 7439 5466
rect 7439 5414 7485 5466
rect 7189 5412 7245 5414
rect 7269 5412 7325 5414
rect 7349 5412 7405 5414
rect 7429 5412 7485 5414
rect 3118 4922 3174 4924
rect 3198 4922 3254 4924
rect 3278 4922 3334 4924
rect 3358 4922 3414 4924
rect 3118 4870 3164 4922
rect 3164 4870 3174 4922
rect 3198 4870 3228 4922
rect 3228 4870 3240 4922
rect 3240 4870 3254 4922
rect 3278 4870 3292 4922
rect 3292 4870 3304 4922
rect 3304 4870 3334 4922
rect 3358 4870 3368 4922
rect 3368 4870 3414 4922
rect 3118 4868 3174 4870
rect 3198 4868 3254 4870
rect 3278 4868 3334 4870
rect 3358 4868 3414 4870
rect 5832 4922 5888 4924
rect 5912 4922 5968 4924
rect 5992 4922 6048 4924
rect 6072 4922 6128 4924
rect 5832 4870 5878 4922
rect 5878 4870 5888 4922
rect 5912 4870 5942 4922
rect 5942 4870 5954 4922
rect 5954 4870 5968 4922
rect 5992 4870 6006 4922
rect 6006 4870 6018 4922
rect 6018 4870 6048 4922
rect 6072 4870 6082 4922
rect 6082 4870 6128 4922
rect 5832 4868 5888 4870
rect 5912 4868 5968 4870
rect 5992 4868 6048 4870
rect 6072 4868 6128 4870
rect 8546 4922 8602 4924
rect 8626 4922 8682 4924
rect 8706 4922 8762 4924
rect 8786 4922 8842 4924
rect 8546 4870 8592 4922
rect 8592 4870 8602 4922
rect 8626 4870 8656 4922
rect 8656 4870 8668 4922
rect 8668 4870 8682 4922
rect 8706 4870 8720 4922
rect 8720 4870 8732 4922
rect 8732 4870 8762 4922
rect 8786 4870 8796 4922
rect 8796 4870 8842 4922
rect 8546 4868 8602 4870
rect 8626 4868 8682 4870
rect 8706 4868 8762 4870
rect 8786 4868 8842 4870
rect 9903 5466 9959 5468
rect 9983 5466 10039 5468
rect 10063 5466 10119 5468
rect 10143 5466 10199 5468
rect 9903 5414 9949 5466
rect 9949 5414 9959 5466
rect 9983 5414 10013 5466
rect 10013 5414 10025 5466
rect 10025 5414 10039 5466
rect 10063 5414 10077 5466
rect 10077 5414 10089 5466
rect 10089 5414 10119 5466
rect 10143 5414 10153 5466
rect 10153 5414 10199 5466
rect 9903 5412 9959 5414
rect 9983 5412 10039 5414
rect 10063 5412 10119 5414
rect 10143 5412 10199 5414
rect 11260 10362 11316 10364
rect 11340 10362 11396 10364
rect 11420 10362 11476 10364
rect 11500 10362 11556 10364
rect 11260 10310 11306 10362
rect 11306 10310 11316 10362
rect 11340 10310 11370 10362
rect 11370 10310 11382 10362
rect 11382 10310 11396 10362
rect 11420 10310 11434 10362
rect 11434 10310 11446 10362
rect 11446 10310 11476 10362
rect 11500 10310 11510 10362
rect 11510 10310 11556 10362
rect 11260 10308 11316 10310
rect 11340 10308 11396 10310
rect 11420 10308 11476 10310
rect 11500 10308 11556 10310
rect 11260 9274 11316 9276
rect 11340 9274 11396 9276
rect 11420 9274 11476 9276
rect 11500 9274 11556 9276
rect 11260 9222 11306 9274
rect 11306 9222 11316 9274
rect 11340 9222 11370 9274
rect 11370 9222 11382 9274
rect 11382 9222 11396 9274
rect 11420 9222 11434 9274
rect 11434 9222 11446 9274
rect 11446 9222 11476 9274
rect 11500 9222 11510 9274
rect 11510 9222 11556 9274
rect 11260 9220 11316 9222
rect 11340 9220 11396 9222
rect 11420 9220 11476 9222
rect 11500 9220 11556 9222
rect 11260 8186 11316 8188
rect 11340 8186 11396 8188
rect 11420 8186 11476 8188
rect 11500 8186 11556 8188
rect 11260 8134 11306 8186
rect 11306 8134 11316 8186
rect 11340 8134 11370 8186
rect 11370 8134 11382 8186
rect 11382 8134 11396 8186
rect 11420 8134 11434 8186
rect 11434 8134 11446 8186
rect 11446 8134 11476 8186
rect 11500 8134 11510 8186
rect 11510 8134 11556 8186
rect 11260 8132 11316 8134
rect 11340 8132 11396 8134
rect 11420 8132 11476 8134
rect 11500 8132 11556 8134
rect 11260 7098 11316 7100
rect 11340 7098 11396 7100
rect 11420 7098 11476 7100
rect 11500 7098 11556 7100
rect 11260 7046 11306 7098
rect 11306 7046 11316 7098
rect 11340 7046 11370 7098
rect 11370 7046 11382 7098
rect 11382 7046 11396 7098
rect 11420 7046 11434 7098
rect 11434 7046 11446 7098
rect 11446 7046 11476 7098
rect 11500 7046 11510 7098
rect 11510 7046 11556 7098
rect 11260 7044 11316 7046
rect 11340 7044 11396 7046
rect 11420 7044 11476 7046
rect 11500 7044 11556 7046
rect 11260 6010 11316 6012
rect 11340 6010 11396 6012
rect 11420 6010 11476 6012
rect 11500 6010 11556 6012
rect 11260 5958 11306 6010
rect 11306 5958 11316 6010
rect 11340 5958 11370 6010
rect 11370 5958 11382 6010
rect 11382 5958 11396 6010
rect 11420 5958 11434 6010
rect 11434 5958 11446 6010
rect 11446 5958 11476 6010
rect 11500 5958 11510 6010
rect 11510 5958 11556 6010
rect 11260 5956 11316 5958
rect 11340 5956 11396 5958
rect 11420 5956 11476 5958
rect 11500 5956 11556 5958
rect 11260 4922 11316 4924
rect 11340 4922 11396 4924
rect 11420 4922 11476 4924
rect 11500 4922 11556 4924
rect 11260 4870 11306 4922
rect 11306 4870 11316 4922
rect 11340 4870 11370 4922
rect 11370 4870 11382 4922
rect 11382 4870 11396 4922
rect 11420 4870 11434 4922
rect 11434 4870 11446 4922
rect 11446 4870 11476 4922
rect 11500 4870 11510 4922
rect 11510 4870 11556 4922
rect 11260 4868 11316 4870
rect 11340 4868 11396 4870
rect 11420 4868 11476 4870
rect 11500 4868 11556 4870
rect 1761 4378 1817 4380
rect 1841 4378 1897 4380
rect 1921 4378 1977 4380
rect 2001 4378 2057 4380
rect 1761 4326 1807 4378
rect 1807 4326 1817 4378
rect 1841 4326 1871 4378
rect 1871 4326 1883 4378
rect 1883 4326 1897 4378
rect 1921 4326 1935 4378
rect 1935 4326 1947 4378
rect 1947 4326 1977 4378
rect 2001 4326 2011 4378
rect 2011 4326 2057 4378
rect 1761 4324 1817 4326
rect 1841 4324 1897 4326
rect 1921 4324 1977 4326
rect 2001 4324 2057 4326
rect 4475 4378 4531 4380
rect 4555 4378 4611 4380
rect 4635 4378 4691 4380
rect 4715 4378 4771 4380
rect 4475 4326 4521 4378
rect 4521 4326 4531 4378
rect 4555 4326 4585 4378
rect 4585 4326 4597 4378
rect 4597 4326 4611 4378
rect 4635 4326 4649 4378
rect 4649 4326 4661 4378
rect 4661 4326 4691 4378
rect 4715 4326 4725 4378
rect 4725 4326 4771 4378
rect 4475 4324 4531 4326
rect 4555 4324 4611 4326
rect 4635 4324 4691 4326
rect 4715 4324 4771 4326
rect 7189 4378 7245 4380
rect 7269 4378 7325 4380
rect 7349 4378 7405 4380
rect 7429 4378 7485 4380
rect 7189 4326 7235 4378
rect 7235 4326 7245 4378
rect 7269 4326 7299 4378
rect 7299 4326 7311 4378
rect 7311 4326 7325 4378
rect 7349 4326 7363 4378
rect 7363 4326 7375 4378
rect 7375 4326 7405 4378
rect 7429 4326 7439 4378
rect 7439 4326 7485 4378
rect 7189 4324 7245 4326
rect 7269 4324 7325 4326
rect 7349 4324 7405 4326
rect 7429 4324 7485 4326
rect 9903 4378 9959 4380
rect 9983 4378 10039 4380
rect 10063 4378 10119 4380
rect 10143 4378 10199 4380
rect 9903 4326 9949 4378
rect 9949 4326 9959 4378
rect 9983 4326 10013 4378
rect 10013 4326 10025 4378
rect 10025 4326 10039 4378
rect 10063 4326 10077 4378
rect 10077 4326 10089 4378
rect 10089 4326 10119 4378
rect 10143 4326 10153 4378
rect 10153 4326 10199 4378
rect 9903 4324 9959 4326
rect 9983 4324 10039 4326
rect 10063 4324 10119 4326
rect 10143 4324 10199 4326
rect 3118 3834 3174 3836
rect 3198 3834 3254 3836
rect 3278 3834 3334 3836
rect 3358 3834 3414 3836
rect 3118 3782 3164 3834
rect 3164 3782 3174 3834
rect 3198 3782 3228 3834
rect 3228 3782 3240 3834
rect 3240 3782 3254 3834
rect 3278 3782 3292 3834
rect 3292 3782 3304 3834
rect 3304 3782 3334 3834
rect 3358 3782 3368 3834
rect 3368 3782 3414 3834
rect 3118 3780 3174 3782
rect 3198 3780 3254 3782
rect 3278 3780 3334 3782
rect 3358 3780 3414 3782
rect 5832 3834 5888 3836
rect 5912 3834 5968 3836
rect 5992 3834 6048 3836
rect 6072 3834 6128 3836
rect 5832 3782 5878 3834
rect 5878 3782 5888 3834
rect 5912 3782 5942 3834
rect 5942 3782 5954 3834
rect 5954 3782 5968 3834
rect 5992 3782 6006 3834
rect 6006 3782 6018 3834
rect 6018 3782 6048 3834
rect 6072 3782 6082 3834
rect 6082 3782 6128 3834
rect 5832 3780 5888 3782
rect 5912 3780 5968 3782
rect 5992 3780 6048 3782
rect 6072 3780 6128 3782
rect 8546 3834 8602 3836
rect 8626 3834 8682 3836
rect 8706 3834 8762 3836
rect 8786 3834 8842 3836
rect 8546 3782 8592 3834
rect 8592 3782 8602 3834
rect 8626 3782 8656 3834
rect 8656 3782 8668 3834
rect 8668 3782 8682 3834
rect 8706 3782 8720 3834
rect 8720 3782 8732 3834
rect 8732 3782 8762 3834
rect 8786 3782 8796 3834
rect 8796 3782 8842 3834
rect 8546 3780 8602 3782
rect 8626 3780 8682 3782
rect 8706 3780 8762 3782
rect 8786 3780 8842 3782
rect 11260 3834 11316 3836
rect 11340 3834 11396 3836
rect 11420 3834 11476 3836
rect 11500 3834 11556 3836
rect 11260 3782 11306 3834
rect 11306 3782 11316 3834
rect 11340 3782 11370 3834
rect 11370 3782 11382 3834
rect 11382 3782 11396 3834
rect 11420 3782 11434 3834
rect 11434 3782 11446 3834
rect 11446 3782 11476 3834
rect 11500 3782 11510 3834
rect 11510 3782 11556 3834
rect 11260 3780 11316 3782
rect 11340 3780 11396 3782
rect 11420 3780 11476 3782
rect 11500 3780 11556 3782
rect 1761 3290 1817 3292
rect 1841 3290 1897 3292
rect 1921 3290 1977 3292
rect 2001 3290 2057 3292
rect 1761 3238 1807 3290
rect 1807 3238 1817 3290
rect 1841 3238 1871 3290
rect 1871 3238 1883 3290
rect 1883 3238 1897 3290
rect 1921 3238 1935 3290
rect 1935 3238 1947 3290
rect 1947 3238 1977 3290
rect 2001 3238 2011 3290
rect 2011 3238 2057 3290
rect 1761 3236 1817 3238
rect 1841 3236 1897 3238
rect 1921 3236 1977 3238
rect 2001 3236 2057 3238
rect 4475 3290 4531 3292
rect 4555 3290 4611 3292
rect 4635 3290 4691 3292
rect 4715 3290 4771 3292
rect 4475 3238 4521 3290
rect 4521 3238 4531 3290
rect 4555 3238 4585 3290
rect 4585 3238 4597 3290
rect 4597 3238 4611 3290
rect 4635 3238 4649 3290
rect 4649 3238 4661 3290
rect 4661 3238 4691 3290
rect 4715 3238 4725 3290
rect 4725 3238 4771 3290
rect 4475 3236 4531 3238
rect 4555 3236 4611 3238
rect 4635 3236 4691 3238
rect 4715 3236 4771 3238
rect 7189 3290 7245 3292
rect 7269 3290 7325 3292
rect 7349 3290 7405 3292
rect 7429 3290 7485 3292
rect 7189 3238 7235 3290
rect 7235 3238 7245 3290
rect 7269 3238 7299 3290
rect 7299 3238 7311 3290
rect 7311 3238 7325 3290
rect 7349 3238 7363 3290
rect 7363 3238 7375 3290
rect 7375 3238 7405 3290
rect 7429 3238 7439 3290
rect 7439 3238 7485 3290
rect 7189 3236 7245 3238
rect 7269 3236 7325 3238
rect 7349 3236 7405 3238
rect 7429 3236 7485 3238
rect 9903 3290 9959 3292
rect 9983 3290 10039 3292
rect 10063 3290 10119 3292
rect 10143 3290 10199 3292
rect 9903 3238 9949 3290
rect 9949 3238 9959 3290
rect 9983 3238 10013 3290
rect 10013 3238 10025 3290
rect 10025 3238 10039 3290
rect 10063 3238 10077 3290
rect 10077 3238 10089 3290
rect 10089 3238 10119 3290
rect 10143 3238 10153 3290
rect 10153 3238 10199 3290
rect 9903 3236 9959 3238
rect 9983 3236 10039 3238
rect 10063 3236 10119 3238
rect 10143 3236 10199 3238
rect 3118 2746 3174 2748
rect 3198 2746 3254 2748
rect 3278 2746 3334 2748
rect 3358 2746 3414 2748
rect 3118 2694 3164 2746
rect 3164 2694 3174 2746
rect 3198 2694 3228 2746
rect 3228 2694 3240 2746
rect 3240 2694 3254 2746
rect 3278 2694 3292 2746
rect 3292 2694 3304 2746
rect 3304 2694 3334 2746
rect 3358 2694 3368 2746
rect 3368 2694 3414 2746
rect 3118 2692 3174 2694
rect 3198 2692 3254 2694
rect 3278 2692 3334 2694
rect 3358 2692 3414 2694
rect 5832 2746 5888 2748
rect 5912 2746 5968 2748
rect 5992 2746 6048 2748
rect 6072 2746 6128 2748
rect 5832 2694 5878 2746
rect 5878 2694 5888 2746
rect 5912 2694 5942 2746
rect 5942 2694 5954 2746
rect 5954 2694 5968 2746
rect 5992 2694 6006 2746
rect 6006 2694 6018 2746
rect 6018 2694 6048 2746
rect 6072 2694 6082 2746
rect 6082 2694 6128 2746
rect 5832 2692 5888 2694
rect 5912 2692 5968 2694
rect 5992 2692 6048 2694
rect 6072 2692 6128 2694
rect 8546 2746 8602 2748
rect 8626 2746 8682 2748
rect 8706 2746 8762 2748
rect 8786 2746 8842 2748
rect 8546 2694 8592 2746
rect 8592 2694 8602 2746
rect 8626 2694 8656 2746
rect 8656 2694 8668 2746
rect 8668 2694 8682 2746
rect 8706 2694 8720 2746
rect 8720 2694 8732 2746
rect 8732 2694 8762 2746
rect 8786 2694 8796 2746
rect 8796 2694 8842 2746
rect 8546 2692 8602 2694
rect 8626 2692 8682 2694
rect 8706 2692 8762 2694
rect 8786 2692 8842 2694
rect 11260 2746 11316 2748
rect 11340 2746 11396 2748
rect 11420 2746 11476 2748
rect 11500 2746 11556 2748
rect 11260 2694 11306 2746
rect 11306 2694 11316 2746
rect 11340 2694 11370 2746
rect 11370 2694 11382 2746
rect 11382 2694 11396 2746
rect 11420 2694 11434 2746
rect 11434 2694 11446 2746
rect 11446 2694 11476 2746
rect 11500 2694 11510 2746
rect 11510 2694 11556 2746
rect 11260 2692 11316 2694
rect 11340 2692 11396 2694
rect 11420 2692 11476 2694
rect 11500 2692 11556 2694
rect 1761 2202 1817 2204
rect 1841 2202 1897 2204
rect 1921 2202 1977 2204
rect 2001 2202 2057 2204
rect 1761 2150 1807 2202
rect 1807 2150 1817 2202
rect 1841 2150 1871 2202
rect 1871 2150 1883 2202
rect 1883 2150 1897 2202
rect 1921 2150 1935 2202
rect 1935 2150 1947 2202
rect 1947 2150 1977 2202
rect 2001 2150 2011 2202
rect 2011 2150 2057 2202
rect 1761 2148 1817 2150
rect 1841 2148 1897 2150
rect 1921 2148 1977 2150
rect 2001 2148 2057 2150
rect 4475 2202 4531 2204
rect 4555 2202 4611 2204
rect 4635 2202 4691 2204
rect 4715 2202 4771 2204
rect 4475 2150 4521 2202
rect 4521 2150 4531 2202
rect 4555 2150 4585 2202
rect 4585 2150 4597 2202
rect 4597 2150 4611 2202
rect 4635 2150 4649 2202
rect 4649 2150 4661 2202
rect 4661 2150 4691 2202
rect 4715 2150 4725 2202
rect 4725 2150 4771 2202
rect 4475 2148 4531 2150
rect 4555 2148 4611 2150
rect 4635 2148 4691 2150
rect 4715 2148 4771 2150
rect 7189 2202 7245 2204
rect 7269 2202 7325 2204
rect 7349 2202 7405 2204
rect 7429 2202 7485 2204
rect 7189 2150 7235 2202
rect 7235 2150 7245 2202
rect 7269 2150 7299 2202
rect 7299 2150 7311 2202
rect 7311 2150 7325 2202
rect 7349 2150 7363 2202
rect 7363 2150 7375 2202
rect 7375 2150 7405 2202
rect 7429 2150 7439 2202
rect 7439 2150 7485 2202
rect 7189 2148 7245 2150
rect 7269 2148 7325 2150
rect 7349 2148 7405 2150
rect 7429 2148 7485 2150
rect 9903 2202 9959 2204
rect 9983 2202 10039 2204
rect 10063 2202 10119 2204
rect 10143 2202 10199 2204
rect 9903 2150 9949 2202
rect 9949 2150 9959 2202
rect 9983 2150 10013 2202
rect 10013 2150 10025 2202
rect 10025 2150 10039 2202
rect 10063 2150 10077 2202
rect 10077 2150 10089 2202
rect 10089 2150 10119 2202
rect 10143 2150 10153 2202
rect 10153 2150 10199 2202
rect 9903 2148 9959 2150
rect 9983 2148 10039 2150
rect 10063 2148 10119 2150
rect 10143 2148 10199 2150
rect 3118 1658 3174 1660
rect 3198 1658 3254 1660
rect 3278 1658 3334 1660
rect 3358 1658 3414 1660
rect 3118 1606 3164 1658
rect 3164 1606 3174 1658
rect 3198 1606 3228 1658
rect 3228 1606 3240 1658
rect 3240 1606 3254 1658
rect 3278 1606 3292 1658
rect 3292 1606 3304 1658
rect 3304 1606 3334 1658
rect 3358 1606 3368 1658
rect 3368 1606 3414 1658
rect 3118 1604 3174 1606
rect 3198 1604 3254 1606
rect 3278 1604 3334 1606
rect 3358 1604 3414 1606
rect 5832 1658 5888 1660
rect 5912 1658 5968 1660
rect 5992 1658 6048 1660
rect 6072 1658 6128 1660
rect 5832 1606 5878 1658
rect 5878 1606 5888 1658
rect 5912 1606 5942 1658
rect 5942 1606 5954 1658
rect 5954 1606 5968 1658
rect 5992 1606 6006 1658
rect 6006 1606 6018 1658
rect 6018 1606 6048 1658
rect 6072 1606 6082 1658
rect 6082 1606 6128 1658
rect 5832 1604 5888 1606
rect 5912 1604 5968 1606
rect 5992 1604 6048 1606
rect 6072 1604 6128 1606
rect 8546 1658 8602 1660
rect 8626 1658 8682 1660
rect 8706 1658 8762 1660
rect 8786 1658 8842 1660
rect 8546 1606 8592 1658
rect 8592 1606 8602 1658
rect 8626 1606 8656 1658
rect 8656 1606 8668 1658
rect 8668 1606 8682 1658
rect 8706 1606 8720 1658
rect 8720 1606 8732 1658
rect 8732 1606 8762 1658
rect 8786 1606 8796 1658
rect 8796 1606 8842 1658
rect 8546 1604 8602 1606
rect 8626 1604 8682 1606
rect 8706 1604 8762 1606
rect 8786 1604 8842 1606
rect 11260 1658 11316 1660
rect 11340 1658 11396 1660
rect 11420 1658 11476 1660
rect 11500 1658 11556 1660
rect 11260 1606 11306 1658
rect 11306 1606 11316 1658
rect 11340 1606 11370 1658
rect 11370 1606 11382 1658
rect 11382 1606 11396 1658
rect 11420 1606 11434 1658
rect 11434 1606 11446 1658
rect 11446 1606 11476 1658
rect 11500 1606 11510 1658
rect 11510 1606 11556 1658
rect 11260 1604 11316 1606
rect 11340 1604 11396 1606
rect 11420 1604 11476 1606
rect 11500 1604 11556 1606
rect 1761 1114 1817 1116
rect 1841 1114 1897 1116
rect 1921 1114 1977 1116
rect 2001 1114 2057 1116
rect 1761 1062 1807 1114
rect 1807 1062 1817 1114
rect 1841 1062 1871 1114
rect 1871 1062 1883 1114
rect 1883 1062 1897 1114
rect 1921 1062 1935 1114
rect 1935 1062 1947 1114
rect 1947 1062 1977 1114
rect 2001 1062 2011 1114
rect 2011 1062 2057 1114
rect 1761 1060 1817 1062
rect 1841 1060 1897 1062
rect 1921 1060 1977 1062
rect 2001 1060 2057 1062
rect 4475 1114 4531 1116
rect 4555 1114 4611 1116
rect 4635 1114 4691 1116
rect 4715 1114 4771 1116
rect 4475 1062 4521 1114
rect 4521 1062 4531 1114
rect 4555 1062 4585 1114
rect 4585 1062 4597 1114
rect 4597 1062 4611 1114
rect 4635 1062 4649 1114
rect 4649 1062 4661 1114
rect 4661 1062 4691 1114
rect 4715 1062 4725 1114
rect 4725 1062 4771 1114
rect 4475 1060 4531 1062
rect 4555 1060 4611 1062
rect 4635 1060 4691 1062
rect 4715 1060 4771 1062
rect 7189 1114 7245 1116
rect 7269 1114 7325 1116
rect 7349 1114 7405 1116
rect 7429 1114 7485 1116
rect 7189 1062 7235 1114
rect 7235 1062 7245 1114
rect 7269 1062 7299 1114
rect 7299 1062 7311 1114
rect 7311 1062 7325 1114
rect 7349 1062 7363 1114
rect 7363 1062 7375 1114
rect 7375 1062 7405 1114
rect 7429 1062 7439 1114
rect 7439 1062 7485 1114
rect 7189 1060 7245 1062
rect 7269 1060 7325 1062
rect 7349 1060 7405 1062
rect 7429 1060 7485 1062
rect 9903 1114 9959 1116
rect 9983 1114 10039 1116
rect 10063 1114 10119 1116
rect 10143 1114 10199 1116
rect 9903 1062 9949 1114
rect 9949 1062 9959 1114
rect 9983 1062 10013 1114
rect 10013 1062 10025 1114
rect 10025 1062 10039 1114
rect 10063 1062 10077 1114
rect 10077 1062 10089 1114
rect 10089 1062 10119 1114
rect 10143 1062 10153 1114
rect 10153 1062 10199 1114
rect 9903 1060 9959 1062
rect 9983 1060 10039 1062
rect 10063 1060 10119 1062
rect 10143 1060 10199 1062
rect 3118 570 3174 572
rect 3198 570 3254 572
rect 3278 570 3334 572
rect 3358 570 3414 572
rect 3118 518 3164 570
rect 3164 518 3174 570
rect 3198 518 3228 570
rect 3228 518 3240 570
rect 3240 518 3254 570
rect 3278 518 3292 570
rect 3292 518 3304 570
rect 3304 518 3334 570
rect 3358 518 3368 570
rect 3368 518 3414 570
rect 3118 516 3174 518
rect 3198 516 3254 518
rect 3278 516 3334 518
rect 3358 516 3414 518
rect 5832 570 5888 572
rect 5912 570 5968 572
rect 5992 570 6048 572
rect 6072 570 6128 572
rect 5832 518 5878 570
rect 5878 518 5888 570
rect 5912 518 5942 570
rect 5942 518 5954 570
rect 5954 518 5968 570
rect 5992 518 6006 570
rect 6006 518 6018 570
rect 6018 518 6048 570
rect 6072 518 6082 570
rect 6082 518 6128 570
rect 5832 516 5888 518
rect 5912 516 5968 518
rect 5992 516 6048 518
rect 6072 516 6128 518
rect 8546 570 8602 572
rect 8626 570 8682 572
rect 8706 570 8762 572
rect 8786 570 8842 572
rect 8546 518 8592 570
rect 8592 518 8602 570
rect 8626 518 8656 570
rect 8656 518 8668 570
rect 8668 518 8682 570
rect 8706 518 8720 570
rect 8720 518 8732 570
rect 8732 518 8762 570
rect 8786 518 8796 570
rect 8796 518 8842 570
rect 8546 516 8602 518
rect 8626 516 8682 518
rect 8706 516 8762 518
rect 8786 516 8842 518
rect 11260 570 11316 572
rect 11340 570 11396 572
rect 11420 570 11476 572
rect 11500 570 11556 572
rect 11260 518 11306 570
rect 11306 518 11316 570
rect 11340 518 11370 570
rect 11370 518 11382 570
rect 11382 518 11396 570
rect 11420 518 11434 570
rect 11434 518 11446 570
rect 11446 518 11476 570
rect 11500 518 11510 570
rect 11510 518 11556 570
rect 11260 516 11316 518
rect 11340 516 11396 518
rect 11420 516 11476 518
rect 11500 516 11556 518
<< metal3 >>
rect 3108 11456 3424 11457
rect 3108 11392 3114 11456
rect 3178 11392 3194 11456
rect 3258 11392 3274 11456
rect 3338 11392 3354 11456
rect 3418 11392 3424 11456
rect 3108 11391 3424 11392
rect 5822 11456 6138 11457
rect 5822 11392 5828 11456
rect 5892 11392 5908 11456
rect 5972 11392 5988 11456
rect 6052 11392 6068 11456
rect 6132 11392 6138 11456
rect 5822 11391 6138 11392
rect 8536 11456 8852 11457
rect 8536 11392 8542 11456
rect 8606 11392 8622 11456
rect 8686 11392 8702 11456
rect 8766 11392 8782 11456
rect 8846 11392 8852 11456
rect 8536 11391 8852 11392
rect 11250 11456 11566 11457
rect 11250 11392 11256 11456
rect 11320 11392 11336 11456
rect 11400 11392 11416 11456
rect 11480 11392 11496 11456
rect 11560 11392 11566 11456
rect 11250 11391 11566 11392
rect 1751 10912 2067 10913
rect 1751 10848 1757 10912
rect 1821 10848 1837 10912
rect 1901 10848 1917 10912
rect 1981 10848 1997 10912
rect 2061 10848 2067 10912
rect 1751 10847 2067 10848
rect 4465 10912 4781 10913
rect 4465 10848 4471 10912
rect 4535 10848 4551 10912
rect 4615 10848 4631 10912
rect 4695 10848 4711 10912
rect 4775 10848 4781 10912
rect 4465 10847 4781 10848
rect 7179 10912 7495 10913
rect 7179 10848 7185 10912
rect 7249 10848 7265 10912
rect 7329 10848 7345 10912
rect 7409 10848 7425 10912
rect 7489 10848 7495 10912
rect 7179 10847 7495 10848
rect 9893 10912 10209 10913
rect 9893 10848 9899 10912
rect 9963 10848 9979 10912
rect 10043 10848 10059 10912
rect 10123 10848 10139 10912
rect 10203 10848 10209 10912
rect 9893 10847 10209 10848
rect 3108 10368 3424 10369
rect 3108 10304 3114 10368
rect 3178 10304 3194 10368
rect 3258 10304 3274 10368
rect 3338 10304 3354 10368
rect 3418 10304 3424 10368
rect 3108 10303 3424 10304
rect 5822 10368 6138 10369
rect 5822 10304 5828 10368
rect 5892 10304 5908 10368
rect 5972 10304 5988 10368
rect 6052 10304 6068 10368
rect 6132 10304 6138 10368
rect 5822 10303 6138 10304
rect 8536 10368 8852 10369
rect 8536 10304 8542 10368
rect 8606 10304 8622 10368
rect 8686 10304 8702 10368
rect 8766 10304 8782 10368
rect 8846 10304 8852 10368
rect 8536 10303 8852 10304
rect 11250 10368 11566 10369
rect 11250 10304 11256 10368
rect 11320 10304 11336 10368
rect 11400 10304 11416 10368
rect 11480 10304 11496 10368
rect 11560 10304 11566 10368
rect 11250 10303 11566 10304
rect 5441 10026 5507 10029
rect 9765 10026 9831 10029
rect 5441 10024 9831 10026
rect 5441 9968 5446 10024
rect 5502 9968 9770 10024
rect 9826 9968 9831 10024
rect 5441 9966 9831 9968
rect 5441 9963 5507 9966
rect 9765 9963 9831 9966
rect 1751 9824 2067 9825
rect 1751 9760 1757 9824
rect 1821 9760 1837 9824
rect 1901 9760 1917 9824
rect 1981 9760 1997 9824
rect 2061 9760 2067 9824
rect 1751 9759 2067 9760
rect 4465 9824 4781 9825
rect 4465 9760 4471 9824
rect 4535 9760 4551 9824
rect 4615 9760 4631 9824
rect 4695 9760 4711 9824
rect 4775 9760 4781 9824
rect 4465 9759 4781 9760
rect 7179 9824 7495 9825
rect 7179 9760 7185 9824
rect 7249 9760 7265 9824
rect 7329 9760 7345 9824
rect 7409 9760 7425 9824
rect 7489 9760 7495 9824
rect 7179 9759 7495 9760
rect 9893 9824 10209 9825
rect 9893 9760 9899 9824
rect 9963 9760 9979 9824
rect 10043 9760 10059 9824
rect 10123 9760 10139 9824
rect 10203 9760 10209 9824
rect 9893 9759 10209 9760
rect 1209 9618 1275 9621
rect 3325 9618 3391 9621
rect 9070 9618 9076 9620
rect 1209 9616 3391 9618
rect 1209 9560 1214 9616
rect 1270 9560 3330 9616
rect 3386 9560 3391 9616
rect 1209 9558 3391 9560
rect 1209 9555 1275 9558
rect 3325 9555 3391 9558
rect 5030 9558 9076 9618
rect 3049 9482 3115 9485
rect 5030 9482 5090 9558
rect 9070 9556 9076 9558
rect 9140 9618 9146 9620
rect 9305 9618 9371 9621
rect 9140 9616 9371 9618
rect 9140 9560 9310 9616
rect 9366 9560 9371 9616
rect 9140 9558 9371 9560
rect 9140 9556 9146 9558
rect 9305 9555 9371 9558
rect 3049 9480 5090 9482
rect 3049 9424 3054 9480
rect 3110 9424 5090 9480
rect 3049 9422 5090 9424
rect 5257 9482 5323 9485
rect 6821 9482 6887 9485
rect 5257 9480 6887 9482
rect 5257 9424 5262 9480
rect 5318 9424 6826 9480
rect 6882 9424 6887 9480
rect 5257 9422 6887 9424
rect 3049 9419 3115 9422
rect 5257 9419 5323 9422
rect 6821 9419 6887 9422
rect 7281 9482 7347 9485
rect 8661 9482 8727 9485
rect 7281 9480 8727 9482
rect 7281 9424 7286 9480
rect 7342 9424 8666 9480
rect 8722 9424 8727 9480
rect 7281 9422 8727 9424
rect 7281 9419 7347 9422
rect 8661 9419 8727 9422
rect 3108 9280 3424 9281
rect 3108 9216 3114 9280
rect 3178 9216 3194 9280
rect 3258 9216 3274 9280
rect 3338 9216 3354 9280
rect 3418 9216 3424 9280
rect 3108 9215 3424 9216
rect 5822 9280 6138 9281
rect 5822 9216 5828 9280
rect 5892 9216 5908 9280
rect 5972 9216 5988 9280
rect 6052 9216 6068 9280
rect 6132 9216 6138 9280
rect 5822 9215 6138 9216
rect 8536 9280 8852 9281
rect 8536 9216 8542 9280
rect 8606 9216 8622 9280
rect 8686 9216 8702 9280
rect 8766 9216 8782 9280
rect 8846 9216 8852 9280
rect 8536 9215 8852 9216
rect 11250 9280 11566 9281
rect 11250 9216 11256 9280
rect 11320 9216 11336 9280
rect 11400 9216 11416 9280
rect 11480 9216 11496 9280
rect 11560 9216 11566 9280
rect 11250 9215 11566 9216
rect 1751 8736 2067 8737
rect 1751 8672 1757 8736
rect 1821 8672 1837 8736
rect 1901 8672 1917 8736
rect 1981 8672 1997 8736
rect 2061 8672 2067 8736
rect 1751 8671 2067 8672
rect 4465 8736 4781 8737
rect 4465 8672 4471 8736
rect 4535 8672 4551 8736
rect 4615 8672 4631 8736
rect 4695 8672 4711 8736
rect 4775 8672 4781 8736
rect 4465 8671 4781 8672
rect 7179 8736 7495 8737
rect 7179 8672 7185 8736
rect 7249 8672 7265 8736
rect 7329 8672 7345 8736
rect 7409 8672 7425 8736
rect 7489 8672 7495 8736
rect 7179 8671 7495 8672
rect 9893 8736 10209 8737
rect 9893 8672 9899 8736
rect 9963 8672 9979 8736
rect 10043 8672 10059 8736
rect 10123 8672 10139 8736
rect 10203 8672 10209 8736
rect 9893 8671 10209 8672
rect 3108 8192 3424 8193
rect 3108 8128 3114 8192
rect 3178 8128 3194 8192
rect 3258 8128 3274 8192
rect 3338 8128 3354 8192
rect 3418 8128 3424 8192
rect 3108 8127 3424 8128
rect 5822 8192 6138 8193
rect 5822 8128 5828 8192
rect 5892 8128 5908 8192
rect 5972 8128 5988 8192
rect 6052 8128 6068 8192
rect 6132 8128 6138 8192
rect 5822 8127 6138 8128
rect 8536 8192 8852 8193
rect 8536 8128 8542 8192
rect 8606 8128 8622 8192
rect 8686 8128 8702 8192
rect 8766 8128 8782 8192
rect 8846 8128 8852 8192
rect 8536 8127 8852 8128
rect 11250 8192 11566 8193
rect 11250 8128 11256 8192
rect 11320 8128 11336 8192
rect 11400 8128 11416 8192
rect 11480 8128 11496 8192
rect 11560 8128 11566 8192
rect 11250 8127 11566 8128
rect 1751 7648 2067 7649
rect 1751 7584 1757 7648
rect 1821 7584 1837 7648
rect 1901 7584 1917 7648
rect 1981 7584 1997 7648
rect 2061 7584 2067 7648
rect 1751 7583 2067 7584
rect 4465 7648 4781 7649
rect 4465 7584 4471 7648
rect 4535 7584 4551 7648
rect 4615 7584 4631 7648
rect 4695 7584 4711 7648
rect 4775 7584 4781 7648
rect 4465 7583 4781 7584
rect 7179 7648 7495 7649
rect 7179 7584 7185 7648
rect 7249 7584 7265 7648
rect 7329 7584 7345 7648
rect 7409 7584 7425 7648
rect 7489 7584 7495 7648
rect 7179 7583 7495 7584
rect 9893 7648 10209 7649
rect 9893 7584 9899 7648
rect 9963 7584 9979 7648
rect 10043 7584 10059 7648
rect 10123 7584 10139 7648
rect 10203 7584 10209 7648
rect 9893 7583 10209 7584
rect 3108 7104 3424 7105
rect 3108 7040 3114 7104
rect 3178 7040 3194 7104
rect 3258 7040 3274 7104
rect 3338 7040 3354 7104
rect 3418 7040 3424 7104
rect 3108 7039 3424 7040
rect 5822 7104 6138 7105
rect 5822 7040 5828 7104
rect 5892 7040 5908 7104
rect 5972 7040 5988 7104
rect 6052 7040 6068 7104
rect 6132 7040 6138 7104
rect 5822 7039 6138 7040
rect 8536 7104 8852 7105
rect 8536 7040 8542 7104
rect 8606 7040 8622 7104
rect 8686 7040 8702 7104
rect 8766 7040 8782 7104
rect 8846 7040 8852 7104
rect 8536 7039 8852 7040
rect 11250 7104 11566 7105
rect 11250 7040 11256 7104
rect 11320 7040 11336 7104
rect 11400 7040 11416 7104
rect 11480 7040 11496 7104
rect 11560 7040 11566 7104
rect 11250 7039 11566 7040
rect 1751 6560 2067 6561
rect 1751 6496 1757 6560
rect 1821 6496 1837 6560
rect 1901 6496 1917 6560
rect 1981 6496 1997 6560
rect 2061 6496 2067 6560
rect 1751 6495 2067 6496
rect 4465 6560 4781 6561
rect 4465 6496 4471 6560
rect 4535 6496 4551 6560
rect 4615 6496 4631 6560
rect 4695 6496 4711 6560
rect 4775 6496 4781 6560
rect 4465 6495 4781 6496
rect 7179 6560 7495 6561
rect 7179 6496 7185 6560
rect 7249 6496 7265 6560
rect 7329 6496 7345 6560
rect 7409 6496 7425 6560
rect 7489 6496 7495 6560
rect 7179 6495 7495 6496
rect 9893 6560 10209 6561
rect 9893 6496 9899 6560
rect 9963 6496 9979 6560
rect 10043 6496 10059 6560
rect 10123 6496 10139 6560
rect 10203 6496 10209 6560
rect 9893 6495 10209 6496
rect 8845 6354 8911 6357
rect 9070 6354 9076 6356
rect 8845 6352 9076 6354
rect 8845 6296 8850 6352
rect 8906 6296 9076 6352
rect 8845 6294 9076 6296
rect 8845 6291 8911 6294
rect 9070 6292 9076 6294
rect 9140 6292 9146 6356
rect 3108 6016 3424 6017
rect 3108 5952 3114 6016
rect 3178 5952 3194 6016
rect 3258 5952 3274 6016
rect 3338 5952 3354 6016
rect 3418 5952 3424 6016
rect 3108 5951 3424 5952
rect 5822 6016 6138 6017
rect 5822 5952 5828 6016
rect 5892 5952 5908 6016
rect 5972 5952 5988 6016
rect 6052 5952 6068 6016
rect 6132 5952 6138 6016
rect 5822 5951 6138 5952
rect 8536 6016 8852 6017
rect 8536 5952 8542 6016
rect 8606 5952 8622 6016
rect 8686 5952 8702 6016
rect 8766 5952 8782 6016
rect 8846 5952 8852 6016
rect 8536 5951 8852 5952
rect 11250 6016 11566 6017
rect 11250 5952 11256 6016
rect 11320 5952 11336 6016
rect 11400 5952 11416 6016
rect 11480 5952 11496 6016
rect 11560 5952 11566 6016
rect 11250 5951 11566 5952
rect 7833 5810 7899 5813
rect 11600 5810 12000 5840
rect 7833 5808 12000 5810
rect 7833 5752 7838 5808
rect 7894 5752 12000 5808
rect 7833 5750 12000 5752
rect 7833 5747 7899 5750
rect 11600 5720 12000 5750
rect 1751 5472 2067 5473
rect 1751 5408 1757 5472
rect 1821 5408 1837 5472
rect 1901 5408 1917 5472
rect 1981 5408 1997 5472
rect 2061 5408 2067 5472
rect 1751 5407 2067 5408
rect 4465 5472 4781 5473
rect 4465 5408 4471 5472
rect 4535 5408 4551 5472
rect 4615 5408 4631 5472
rect 4695 5408 4711 5472
rect 4775 5408 4781 5472
rect 4465 5407 4781 5408
rect 7179 5472 7495 5473
rect 7179 5408 7185 5472
rect 7249 5408 7265 5472
rect 7329 5408 7345 5472
rect 7409 5408 7425 5472
rect 7489 5408 7495 5472
rect 7179 5407 7495 5408
rect 9893 5472 10209 5473
rect 9893 5408 9899 5472
rect 9963 5408 9979 5472
rect 10043 5408 10059 5472
rect 10123 5408 10139 5472
rect 10203 5408 10209 5472
rect 9893 5407 10209 5408
rect 3108 4928 3424 4929
rect 3108 4864 3114 4928
rect 3178 4864 3194 4928
rect 3258 4864 3274 4928
rect 3338 4864 3354 4928
rect 3418 4864 3424 4928
rect 3108 4863 3424 4864
rect 5822 4928 6138 4929
rect 5822 4864 5828 4928
rect 5892 4864 5908 4928
rect 5972 4864 5988 4928
rect 6052 4864 6068 4928
rect 6132 4864 6138 4928
rect 5822 4863 6138 4864
rect 8536 4928 8852 4929
rect 8536 4864 8542 4928
rect 8606 4864 8622 4928
rect 8686 4864 8702 4928
rect 8766 4864 8782 4928
rect 8846 4864 8852 4928
rect 8536 4863 8852 4864
rect 11250 4928 11566 4929
rect 11250 4864 11256 4928
rect 11320 4864 11336 4928
rect 11400 4864 11416 4928
rect 11480 4864 11496 4928
rect 11560 4864 11566 4928
rect 11250 4863 11566 4864
rect 1751 4384 2067 4385
rect 1751 4320 1757 4384
rect 1821 4320 1837 4384
rect 1901 4320 1917 4384
rect 1981 4320 1997 4384
rect 2061 4320 2067 4384
rect 1751 4319 2067 4320
rect 4465 4384 4781 4385
rect 4465 4320 4471 4384
rect 4535 4320 4551 4384
rect 4615 4320 4631 4384
rect 4695 4320 4711 4384
rect 4775 4320 4781 4384
rect 4465 4319 4781 4320
rect 7179 4384 7495 4385
rect 7179 4320 7185 4384
rect 7249 4320 7265 4384
rect 7329 4320 7345 4384
rect 7409 4320 7425 4384
rect 7489 4320 7495 4384
rect 7179 4319 7495 4320
rect 9893 4384 10209 4385
rect 9893 4320 9899 4384
rect 9963 4320 9979 4384
rect 10043 4320 10059 4384
rect 10123 4320 10139 4384
rect 10203 4320 10209 4384
rect 9893 4319 10209 4320
rect 3108 3840 3424 3841
rect 3108 3776 3114 3840
rect 3178 3776 3194 3840
rect 3258 3776 3274 3840
rect 3338 3776 3354 3840
rect 3418 3776 3424 3840
rect 3108 3775 3424 3776
rect 5822 3840 6138 3841
rect 5822 3776 5828 3840
rect 5892 3776 5908 3840
rect 5972 3776 5988 3840
rect 6052 3776 6068 3840
rect 6132 3776 6138 3840
rect 5822 3775 6138 3776
rect 8536 3840 8852 3841
rect 8536 3776 8542 3840
rect 8606 3776 8622 3840
rect 8686 3776 8702 3840
rect 8766 3776 8782 3840
rect 8846 3776 8852 3840
rect 8536 3775 8852 3776
rect 11250 3840 11566 3841
rect 11250 3776 11256 3840
rect 11320 3776 11336 3840
rect 11400 3776 11416 3840
rect 11480 3776 11496 3840
rect 11560 3776 11566 3840
rect 11250 3775 11566 3776
rect 1751 3296 2067 3297
rect 1751 3232 1757 3296
rect 1821 3232 1837 3296
rect 1901 3232 1917 3296
rect 1981 3232 1997 3296
rect 2061 3232 2067 3296
rect 1751 3231 2067 3232
rect 4465 3296 4781 3297
rect 4465 3232 4471 3296
rect 4535 3232 4551 3296
rect 4615 3232 4631 3296
rect 4695 3232 4711 3296
rect 4775 3232 4781 3296
rect 4465 3231 4781 3232
rect 7179 3296 7495 3297
rect 7179 3232 7185 3296
rect 7249 3232 7265 3296
rect 7329 3232 7345 3296
rect 7409 3232 7425 3296
rect 7489 3232 7495 3296
rect 7179 3231 7495 3232
rect 9893 3296 10209 3297
rect 9893 3232 9899 3296
rect 9963 3232 9979 3296
rect 10043 3232 10059 3296
rect 10123 3232 10139 3296
rect 10203 3232 10209 3296
rect 9893 3231 10209 3232
rect 3108 2752 3424 2753
rect 3108 2688 3114 2752
rect 3178 2688 3194 2752
rect 3258 2688 3274 2752
rect 3338 2688 3354 2752
rect 3418 2688 3424 2752
rect 3108 2687 3424 2688
rect 5822 2752 6138 2753
rect 5822 2688 5828 2752
rect 5892 2688 5908 2752
rect 5972 2688 5988 2752
rect 6052 2688 6068 2752
rect 6132 2688 6138 2752
rect 5822 2687 6138 2688
rect 8536 2752 8852 2753
rect 8536 2688 8542 2752
rect 8606 2688 8622 2752
rect 8686 2688 8702 2752
rect 8766 2688 8782 2752
rect 8846 2688 8852 2752
rect 8536 2687 8852 2688
rect 11250 2752 11566 2753
rect 11250 2688 11256 2752
rect 11320 2688 11336 2752
rect 11400 2688 11416 2752
rect 11480 2688 11496 2752
rect 11560 2688 11566 2752
rect 11250 2687 11566 2688
rect 1751 2208 2067 2209
rect 1751 2144 1757 2208
rect 1821 2144 1837 2208
rect 1901 2144 1917 2208
rect 1981 2144 1997 2208
rect 2061 2144 2067 2208
rect 1751 2143 2067 2144
rect 4465 2208 4781 2209
rect 4465 2144 4471 2208
rect 4535 2144 4551 2208
rect 4615 2144 4631 2208
rect 4695 2144 4711 2208
rect 4775 2144 4781 2208
rect 4465 2143 4781 2144
rect 7179 2208 7495 2209
rect 7179 2144 7185 2208
rect 7249 2144 7265 2208
rect 7329 2144 7345 2208
rect 7409 2144 7425 2208
rect 7489 2144 7495 2208
rect 7179 2143 7495 2144
rect 9893 2208 10209 2209
rect 9893 2144 9899 2208
rect 9963 2144 9979 2208
rect 10043 2144 10059 2208
rect 10123 2144 10139 2208
rect 10203 2144 10209 2208
rect 9893 2143 10209 2144
rect 3108 1664 3424 1665
rect 3108 1600 3114 1664
rect 3178 1600 3194 1664
rect 3258 1600 3274 1664
rect 3338 1600 3354 1664
rect 3418 1600 3424 1664
rect 3108 1599 3424 1600
rect 5822 1664 6138 1665
rect 5822 1600 5828 1664
rect 5892 1600 5908 1664
rect 5972 1600 5988 1664
rect 6052 1600 6068 1664
rect 6132 1600 6138 1664
rect 5822 1599 6138 1600
rect 8536 1664 8852 1665
rect 8536 1600 8542 1664
rect 8606 1600 8622 1664
rect 8686 1600 8702 1664
rect 8766 1600 8782 1664
rect 8846 1600 8852 1664
rect 8536 1599 8852 1600
rect 11250 1664 11566 1665
rect 11250 1600 11256 1664
rect 11320 1600 11336 1664
rect 11400 1600 11416 1664
rect 11480 1600 11496 1664
rect 11560 1600 11566 1664
rect 11250 1599 11566 1600
rect 1751 1120 2067 1121
rect 1751 1056 1757 1120
rect 1821 1056 1837 1120
rect 1901 1056 1917 1120
rect 1981 1056 1997 1120
rect 2061 1056 2067 1120
rect 1751 1055 2067 1056
rect 4465 1120 4781 1121
rect 4465 1056 4471 1120
rect 4535 1056 4551 1120
rect 4615 1056 4631 1120
rect 4695 1056 4711 1120
rect 4775 1056 4781 1120
rect 4465 1055 4781 1056
rect 7179 1120 7495 1121
rect 7179 1056 7185 1120
rect 7249 1056 7265 1120
rect 7329 1056 7345 1120
rect 7409 1056 7425 1120
rect 7489 1056 7495 1120
rect 7179 1055 7495 1056
rect 9893 1120 10209 1121
rect 9893 1056 9899 1120
rect 9963 1056 9979 1120
rect 10043 1056 10059 1120
rect 10123 1056 10139 1120
rect 10203 1056 10209 1120
rect 9893 1055 10209 1056
rect 3108 576 3424 577
rect 3108 512 3114 576
rect 3178 512 3194 576
rect 3258 512 3274 576
rect 3338 512 3354 576
rect 3418 512 3424 576
rect 3108 511 3424 512
rect 5822 576 6138 577
rect 5822 512 5828 576
rect 5892 512 5908 576
rect 5972 512 5988 576
rect 6052 512 6068 576
rect 6132 512 6138 576
rect 5822 511 6138 512
rect 8536 576 8852 577
rect 8536 512 8542 576
rect 8606 512 8622 576
rect 8686 512 8702 576
rect 8766 512 8782 576
rect 8846 512 8852 576
rect 8536 511 8852 512
rect 11250 576 11566 577
rect 11250 512 11256 576
rect 11320 512 11336 576
rect 11400 512 11416 576
rect 11480 512 11496 576
rect 11560 512 11566 576
rect 11250 511 11566 512
<< via3 >>
rect 3114 11452 3178 11456
rect 3114 11396 3118 11452
rect 3118 11396 3174 11452
rect 3174 11396 3178 11452
rect 3114 11392 3178 11396
rect 3194 11452 3258 11456
rect 3194 11396 3198 11452
rect 3198 11396 3254 11452
rect 3254 11396 3258 11452
rect 3194 11392 3258 11396
rect 3274 11452 3338 11456
rect 3274 11396 3278 11452
rect 3278 11396 3334 11452
rect 3334 11396 3338 11452
rect 3274 11392 3338 11396
rect 3354 11452 3418 11456
rect 3354 11396 3358 11452
rect 3358 11396 3414 11452
rect 3414 11396 3418 11452
rect 3354 11392 3418 11396
rect 5828 11452 5892 11456
rect 5828 11396 5832 11452
rect 5832 11396 5888 11452
rect 5888 11396 5892 11452
rect 5828 11392 5892 11396
rect 5908 11452 5972 11456
rect 5908 11396 5912 11452
rect 5912 11396 5968 11452
rect 5968 11396 5972 11452
rect 5908 11392 5972 11396
rect 5988 11452 6052 11456
rect 5988 11396 5992 11452
rect 5992 11396 6048 11452
rect 6048 11396 6052 11452
rect 5988 11392 6052 11396
rect 6068 11452 6132 11456
rect 6068 11396 6072 11452
rect 6072 11396 6128 11452
rect 6128 11396 6132 11452
rect 6068 11392 6132 11396
rect 8542 11452 8606 11456
rect 8542 11396 8546 11452
rect 8546 11396 8602 11452
rect 8602 11396 8606 11452
rect 8542 11392 8606 11396
rect 8622 11452 8686 11456
rect 8622 11396 8626 11452
rect 8626 11396 8682 11452
rect 8682 11396 8686 11452
rect 8622 11392 8686 11396
rect 8702 11452 8766 11456
rect 8702 11396 8706 11452
rect 8706 11396 8762 11452
rect 8762 11396 8766 11452
rect 8702 11392 8766 11396
rect 8782 11452 8846 11456
rect 8782 11396 8786 11452
rect 8786 11396 8842 11452
rect 8842 11396 8846 11452
rect 8782 11392 8846 11396
rect 11256 11452 11320 11456
rect 11256 11396 11260 11452
rect 11260 11396 11316 11452
rect 11316 11396 11320 11452
rect 11256 11392 11320 11396
rect 11336 11452 11400 11456
rect 11336 11396 11340 11452
rect 11340 11396 11396 11452
rect 11396 11396 11400 11452
rect 11336 11392 11400 11396
rect 11416 11452 11480 11456
rect 11416 11396 11420 11452
rect 11420 11396 11476 11452
rect 11476 11396 11480 11452
rect 11416 11392 11480 11396
rect 11496 11452 11560 11456
rect 11496 11396 11500 11452
rect 11500 11396 11556 11452
rect 11556 11396 11560 11452
rect 11496 11392 11560 11396
rect 1757 10908 1821 10912
rect 1757 10852 1761 10908
rect 1761 10852 1817 10908
rect 1817 10852 1821 10908
rect 1757 10848 1821 10852
rect 1837 10908 1901 10912
rect 1837 10852 1841 10908
rect 1841 10852 1897 10908
rect 1897 10852 1901 10908
rect 1837 10848 1901 10852
rect 1917 10908 1981 10912
rect 1917 10852 1921 10908
rect 1921 10852 1977 10908
rect 1977 10852 1981 10908
rect 1917 10848 1981 10852
rect 1997 10908 2061 10912
rect 1997 10852 2001 10908
rect 2001 10852 2057 10908
rect 2057 10852 2061 10908
rect 1997 10848 2061 10852
rect 4471 10908 4535 10912
rect 4471 10852 4475 10908
rect 4475 10852 4531 10908
rect 4531 10852 4535 10908
rect 4471 10848 4535 10852
rect 4551 10908 4615 10912
rect 4551 10852 4555 10908
rect 4555 10852 4611 10908
rect 4611 10852 4615 10908
rect 4551 10848 4615 10852
rect 4631 10908 4695 10912
rect 4631 10852 4635 10908
rect 4635 10852 4691 10908
rect 4691 10852 4695 10908
rect 4631 10848 4695 10852
rect 4711 10908 4775 10912
rect 4711 10852 4715 10908
rect 4715 10852 4771 10908
rect 4771 10852 4775 10908
rect 4711 10848 4775 10852
rect 7185 10908 7249 10912
rect 7185 10852 7189 10908
rect 7189 10852 7245 10908
rect 7245 10852 7249 10908
rect 7185 10848 7249 10852
rect 7265 10908 7329 10912
rect 7265 10852 7269 10908
rect 7269 10852 7325 10908
rect 7325 10852 7329 10908
rect 7265 10848 7329 10852
rect 7345 10908 7409 10912
rect 7345 10852 7349 10908
rect 7349 10852 7405 10908
rect 7405 10852 7409 10908
rect 7345 10848 7409 10852
rect 7425 10908 7489 10912
rect 7425 10852 7429 10908
rect 7429 10852 7485 10908
rect 7485 10852 7489 10908
rect 7425 10848 7489 10852
rect 9899 10908 9963 10912
rect 9899 10852 9903 10908
rect 9903 10852 9959 10908
rect 9959 10852 9963 10908
rect 9899 10848 9963 10852
rect 9979 10908 10043 10912
rect 9979 10852 9983 10908
rect 9983 10852 10039 10908
rect 10039 10852 10043 10908
rect 9979 10848 10043 10852
rect 10059 10908 10123 10912
rect 10059 10852 10063 10908
rect 10063 10852 10119 10908
rect 10119 10852 10123 10908
rect 10059 10848 10123 10852
rect 10139 10908 10203 10912
rect 10139 10852 10143 10908
rect 10143 10852 10199 10908
rect 10199 10852 10203 10908
rect 10139 10848 10203 10852
rect 3114 10364 3178 10368
rect 3114 10308 3118 10364
rect 3118 10308 3174 10364
rect 3174 10308 3178 10364
rect 3114 10304 3178 10308
rect 3194 10364 3258 10368
rect 3194 10308 3198 10364
rect 3198 10308 3254 10364
rect 3254 10308 3258 10364
rect 3194 10304 3258 10308
rect 3274 10364 3338 10368
rect 3274 10308 3278 10364
rect 3278 10308 3334 10364
rect 3334 10308 3338 10364
rect 3274 10304 3338 10308
rect 3354 10364 3418 10368
rect 3354 10308 3358 10364
rect 3358 10308 3414 10364
rect 3414 10308 3418 10364
rect 3354 10304 3418 10308
rect 5828 10364 5892 10368
rect 5828 10308 5832 10364
rect 5832 10308 5888 10364
rect 5888 10308 5892 10364
rect 5828 10304 5892 10308
rect 5908 10364 5972 10368
rect 5908 10308 5912 10364
rect 5912 10308 5968 10364
rect 5968 10308 5972 10364
rect 5908 10304 5972 10308
rect 5988 10364 6052 10368
rect 5988 10308 5992 10364
rect 5992 10308 6048 10364
rect 6048 10308 6052 10364
rect 5988 10304 6052 10308
rect 6068 10364 6132 10368
rect 6068 10308 6072 10364
rect 6072 10308 6128 10364
rect 6128 10308 6132 10364
rect 6068 10304 6132 10308
rect 8542 10364 8606 10368
rect 8542 10308 8546 10364
rect 8546 10308 8602 10364
rect 8602 10308 8606 10364
rect 8542 10304 8606 10308
rect 8622 10364 8686 10368
rect 8622 10308 8626 10364
rect 8626 10308 8682 10364
rect 8682 10308 8686 10364
rect 8622 10304 8686 10308
rect 8702 10364 8766 10368
rect 8702 10308 8706 10364
rect 8706 10308 8762 10364
rect 8762 10308 8766 10364
rect 8702 10304 8766 10308
rect 8782 10364 8846 10368
rect 8782 10308 8786 10364
rect 8786 10308 8842 10364
rect 8842 10308 8846 10364
rect 8782 10304 8846 10308
rect 11256 10364 11320 10368
rect 11256 10308 11260 10364
rect 11260 10308 11316 10364
rect 11316 10308 11320 10364
rect 11256 10304 11320 10308
rect 11336 10364 11400 10368
rect 11336 10308 11340 10364
rect 11340 10308 11396 10364
rect 11396 10308 11400 10364
rect 11336 10304 11400 10308
rect 11416 10364 11480 10368
rect 11416 10308 11420 10364
rect 11420 10308 11476 10364
rect 11476 10308 11480 10364
rect 11416 10304 11480 10308
rect 11496 10364 11560 10368
rect 11496 10308 11500 10364
rect 11500 10308 11556 10364
rect 11556 10308 11560 10364
rect 11496 10304 11560 10308
rect 1757 9820 1821 9824
rect 1757 9764 1761 9820
rect 1761 9764 1817 9820
rect 1817 9764 1821 9820
rect 1757 9760 1821 9764
rect 1837 9820 1901 9824
rect 1837 9764 1841 9820
rect 1841 9764 1897 9820
rect 1897 9764 1901 9820
rect 1837 9760 1901 9764
rect 1917 9820 1981 9824
rect 1917 9764 1921 9820
rect 1921 9764 1977 9820
rect 1977 9764 1981 9820
rect 1917 9760 1981 9764
rect 1997 9820 2061 9824
rect 1997 9764 2001 9820
rect 2001 9764 2057 9820
rect 2057 9764 2061 9820
rect 1997 9760 2061 9764
rect 4471 9820 4535 9824
rect 4471 9764 4475 9820
rect 4475 9764 4531 9820
rect 4531 9764 4535 9820
rect 4471 9760 4535 9764
rect 4551 9820 4615 9824
rect 4551 9764 4555 9820
rect 4555 9764 4611 9820
rect 4611 9764 4615 9820
rect 4551 9760 4615 9764
rect 4631 9820 4695 9824
rect 4631 9764 4635 9820
rect 4635 9764 4691 9820
rect 4691 9764 4695 9820
rect 4631 9760 4695 9764
rect 4711 9820 4775 9824
rect 4711 9764 4715 9820
rect 4715 9764 4771 9820
rect 4771 9764 4775 9820
rect 4711 9760 4775 9764
rect 7185 9820 7249 9824
rect 7185 9764 7189 9820
rect 7189 9764 7245 9820
rect 7245 9764 7249 9820
rect 7185 9760 7249 9764
rect 7265 9820 7329 9824
rect 7265 9764 7269 9820
rect 7269 9764 7325 9820
rect 7325 9764 7329 9820
rect 7265 9760 7329 9764
rect 7345 9820 7409 9824
rect 7345 9764 7349 9820
rect 7349 9764 7405 9820
rect 7405 9764 7409 9820
rect 7345 9760 7409 9764
rect 7425 9820 7489 9824
rect 7425 9764 7429 9820
rect 7429 9764 7485 9820
rect 7485 9764 7489 9820
rect 7425 9760 7489 9764
rect 9899 9820 9963 9824
rect 9899 9764 9903 9820
rect 9903 9764 9959 9820
rect 9959 9764 9963 9820
rect 9899 9760 9963 9764
rect 9979 9820 10043 9824
rect 9979 9764 9983 9820
rect 9983 9764 10039 9820
rect 10039 9764 10043 9820
rect 9979 9760 10043 9764
rect 10059 9820 10123 9824
rect 10059 9764 10063 9820
rect 10063 9764 10119 9820
rect 10119 9764 10123 9820
rect 10059 9760 10123 9764
rect 10139 9820 10203 9824
rect 10139 9764 10143 9820
rect 10143 9764 10199 9820
rect 10199 9764 10203 9820
rect 10139 9760 10203 9764
rect 9076 9556 9140 9620
rect 3114 9276 3178 9280
rect 3114 9220 3118 9276
rect 3118 9220 3174 9276
rect 3174 9220 3178 9276
rect 3114 9216 3178 9220
rect 3194 9276 3258 9280
rect 3194 9220 3198 9276
rect 3198 9220 3254 9276
rect 3254 9220 3258 9276
rect 3194 9216 3258 9220
rect 3274 9276 3338 9280
rect 3274 9220 3278 9276
rect 3278 9220 3334 9276
rect 3334 9220 3338 9276
rect 3274 9216 3338 9220
rect 3354 9276 3418 9280
rect 3354 9220 3358 9276
rect 3358 9220 3414 9276
rect 3414 9220 3418 9276
rect 3354 9216 3418 9220
rect 5828 9276 5892 9280
rect 5828 9220 5832 9276
rect 5832 9220 5888 9276
rect 5888 9220 5892 9276
rect 5828 9216 5892 9220
rect 5908 9276 5972 9280
rect 5908 9220 5912 9276
rect 5912 9220 5968 9276
rect 5968 9220 5972 9276
rect 5908 9216 5972 9220
rect 5988 9276 6052 9280
rect 5988 9220 5992 9276
rect 5992 9220 6048 9276
rect 6048 9220 6052 9276
rect 5988 9216 6052 9220
rect 6068 9276 6132 9280
rect 6068 9220 6072 9276
rect 6072 9220 6128 9276
rect 6128 9220 6132 9276
rect 6068 9216 6132 9220
rect 8542 9276 8606 9280
rect 8542 9220 8546 9276
rect 8546 9220 8602 9276
rect 8602 9220 8606 9276
rect 8542 9216 8606 9220
rect 8622 9276 8686 9280
rect 8622 9220 8626 9276
rect 8626 9220 8682 9276
rect 8682 9220 8686 9276
rect 8622 9216 8686 9220
rect 8702 9276 8766 9280
rect 8702 9220 8706 9276
rect 8706 9220 8762 9276
rect 8762 9220 8766 9276
rect 8702 9216 8766 9220
rect 8782 9276 8846 9280
rect 8782 9220 8786 9276
rect 8786 9220 8842 9276
rect 8842 9220 8846 9276
rect 8782 9216 8846 9220
rect 11256 9276 11320 9280
rect 11256 9220 11260 9276
rect 11260 9220 11316 9276
rect 11316 9220 11320 9276
rect 11256 9216 11320 9220
rect 11336 9276 11400 9280
rect 11336 9220 11340 9276
rect 11340 9220 11396 9276
rect 11396 9220 11400 9276
rect 11336 9216 11400 9220
rect 11416 9276 11480 9280
rect 11416 9220 11420 9276
rect 11420 9220 11476 9276
rect 11476 9220 11480 9276
rect 11416 9216 11480 9220
rect 11496 9276 11560 9280
rect 11496 9220 11500 9276
rect 11500 9220 11556 9276
rect 11556 9220 11560 9276
rect 11496 9216 11560 9220
rect 1757 8732 1821 8736
rect 1757 8676 1761 8732
rect 1761 8676 1817 8732
rect 1817 8676 1821 8732
rect 1757 8672 1821 8676
rect 1837 8732 1901 8736
rect 1837 8676 1841 8732
rect 1841 8676 1897 8732
rect 1897 8676 1901 8732
rect 1837 8672 1901 8676
rect 1917 8732 1981 8736
rect 1917 8676 1921 8732
rect 1921 8676 1977 8732
rect 1977 8676 1981 8732
rect 1917 8672 1981 8676
rect 1997 8732 2061 8736
rect 1997 8676 2001 8732
rect 2001 8676 2057 8732
rect 2057 8676 2061 8732
rect 1997 8672 2061 8676
rect 4471 8732 4535 8736
rect 4471 8676 4475 8732
rect 4475 8676 4531 8732
rect 4531 8676 4535 8732
rect 4471 8672 4535 8676
rect 4551 8732 4615 8736
rect 4551 8676 4555 8732
rect 4555 8676 4611 8732
rect 4611 8676 4615 8732
rect 4551 8672 4615 8676
rect 4631 8732 4695 8736
rect 4631 8676 4635 8732
rect 4635 8676 4691 8732
rect 4691 8676 4695 8732
rect 4631 8672 4695 8676
rect 4711 8732 4775 8736
rect 4711 8676 4715 8732
rect 4715 8676 4771 8732
rect 4771 8676 4775 8732
rect 4711 8672 4775 8676
rect 7185 8732 7249 8736
rect 7185 8676 7189 8732
rect 7189 8676 7245 8732
rect 7245 8676 7249 8732
rect 7185 8672 7249 8676
rect 7265 8732 7329 8736
rect 7265 8676 7269 8732
rect 7269 8676 7325 8732
rect 7325 8676 7329 8732
rect 7265 8672 7329 8676
rect 7345 8732 7409 8736
rect 7345 8676 7349 8732
rect 7349 8676 7405 8732
rect 7405 8676 7409 8732
rect 7345 8672 7409 8676
rect 7425 8732 7489 8736
rect 7425 8676 7429 8732
rect 7429 8676 7485 8732
rect 7485 8676 7489 8732
rect 7425 8672 7489 8676
rect 9899 8732 9963 8736
rect 9899 8676 9903 8732
rect 9903 8676 9959 8732
rect 9959 8676 9963 8732
rect 9899 8672 9963 8676
rect 9979 8732 10043 8736
rect 9979 8676 9983 8732
rect 9983 8676 10039 8732
rect 10039 8676 10043 8732
rect 9979 8672 10043 8676
rect 10059 8732 10123 8736
rect 10059 8676 10063 8732
rect 10063 8676 10119 8732
rect 10119 8676 10123 8732
rect 10059 8672 10123 8676
rect 10139 8732 10203 8736
rect 10139 8676 10143 8732
rect 10143 8676 10199 8732
rect 10199 8676 10203 8732
rect 10139 8672 10203 8676
rect 3114 8188 3178 8192
rect 3114 8132 3118 8188
rect 3118 8132 3174 8188
rect 3174 8132 3178 8188
rect 3114 8128 3178 8132
rect 3194 8188 3258 8192
rect 3194 8132 3198 8188
rect 3198 8132 3254 8188
rect 3254 8132 3258 8188
rect 3194 8128 3258 8132
rect 3274 8188 3338 8192
rect 3274 8132 3278 8188
rect 3278 8132 3334 8188
rect 3334 8132 3338 8188
rect 3274 8128 3338 8132
rect 3354 8188 3418 8192
rect 3354 8132 3358 8188
rect 3358 8132 3414 8188
rect 3414 8132 3418 8188
rect 3354 8128 3418 8132
rect 5828 8188 5892 8192
rect 5828 8132 5832 8188
rect 5832 8132 5888 8188
rect 5888 8132 5892 8188
rect 5828 8128 5892 8132
rect 5908 8188 5972 8192
rect 5908 8132 5912 8188
rect 5912 8132 5968 8188
rect 5968 8132 5972 8188
rect 5908 8128 5972 8132
rect 5988 8188 6052 8192
rect 5988 8132 5992 8188
rect 5992 8132 6048 8188
rect 6048 8132 6052 8188
rect 5988 8128 6052 8132
rect 6068 8188 6132 8192
rect 6068 8132 6072 8188
rect 6072 8132 6128 8188
rect 6128 8132 6132 8188
rect 6068 8128 6132 8132
rect 8542 8188 8606 8192
rect 8542 8132 8546 8188
rect 8546 8132 8602 8188
rect 8602 8132 8606 8188
rect 8542 8128 8606 8132
rect 8622 8188 8686 8192
rect 8622 8132 8626 8188
rect 8626 8132 8682 8188
rect 8682 8132 8686 8188
rect 8622 8128 8686 8132
rect 8702 8188 8766 8192
rect 8702 8132 8706 8188
rect 8706 8132 8762 8188
rect 8762 8132 8766 8188
rect 8702 8128 8766 8132
rect 8782 8188 8846 8192
rect 8782 8132 8786 8188
rect 8786 8132 8842 8188
rect 8842 8132 8846 8188
rect 8782 8128 8846 8132
rect 11256 8188 11320 8192
rect 11256 8132 11260 8188
rect 11260 8132 11316 8188
rect 11316 8132 11320 8188
rect 11256 8128 11320 8132
rect 11336 8188 11400 8192
rect 11336 8132 11340 8188
rect 11340 8132 11396 8188
rect 11396 8132 11400 8188
rect 11336 8128 11400 8132
rect 11416 8188 11480 8192
rect 11416 8132 11420 8188
rect 11420 8132 11476 8188
rect 11476 8132 11480 8188
rect 11416 8128 11480 8132
rect 11496 8188 11560 8192
rect 11496 8132 11500 8188
rect 11500 8132 11556 8188
rect 11556 8132 11560 8188
rect 11496 8128 11560 8132
rect 1757 7644 1821 7648
rect 1757 7588 1761 7644
rect 1761 7588 1817 7644
rect 1817 7588 1821 7644
rect 1757 7584 1821 7588
rect 1837 7644 1901 7648
rect 1837 7588 1841 7644
rect 1841 7588 1897 7644
rect 1897 7588 1901 7644
rect 1837 7584 1901 7588
rect 1917 7644 1981 7648
rect 1917 7588 1921 7644
rect 1921 7588 1977 7644
rect 1977 7588 1981 7644
rect 1917 7584 1981 7588
rect 1997 7644 2061 7648
rect 1997 7588 2001 7644
rect 2001 7588 2057 7644
rect 2057 7588 2061 7644
rect 1997 7584 2061 7588
rect 4471 7644 4535 7648
rect 4471 7588 4475 7644
rect 4475 7588 4531 7644
rect 4531 7588 4535 7644
rect 4471 7584 4535 7588
rect 4551 7644 4615 7648
rect 4551 7588 4555 7644
rect 4555 7588 4611 7644
rect 4611 7588 4615 7644
rect 4551 7584 4615 7588
rect 4631 7644 4695 7648
rect 4631 7588 4635 7644
rect 4635 7588 4691 7644
rect 4691 7588 4695 7644
rect 4631 7584 4695 7588
rect 4711 7644 4775 7648
rect 4711 7588 4715 7644
rect 4715 7588 4771 7644
rect 4771 7588 4775 7644
rect 4711 7584 4775 7588
rect 7185 7644 7249 7648
rect 7185 7588 7189 7644
rect 7189 7588 7245 7644
rect 7245 7588 7249 7644
rect 7185 7584 7249 7588
rect 7265 7644 7329 7648
rect 7265 7588 7269 7644
rect 7269 7588 7325 7644
rect 7325 7588 7329 7644
rect 7265 7584 7329 7588
rect 7345 7644 7409 7648
rect 7345 7588 7349 7644
rect 7349 7588 7405 7644
rect 7405 7588 7409 7644
rect 7345 7584 7409 7588
rect 7425 7644 7489 7648
rect 7425 7588 7429 7644
rect 7429 7588 7485 7644
rect 7485 7588 7489 7644
rect 7425 7584 7489 7588
rect 9899 7644 9963 7648
rect 9899 7588 9903 7644
rect 9903 7588 9959 7644
rect 9959 7588 9963 7644
rect 9899 7584 9963 7588
rect 9979 7644 10043 7648
rect 9979 7588 9983 7644
rect 9983 7588 10039 7644
rect 10039 7588 10043 7644
rect 9979 7584 10043 7588
rect 10059 7644 10123 7648
rect 10059 7588 10063 7644
rect 10063 7588 10119 7644
rect 10119 7588 10123 7644
rect 10059 7584 10123 7588
rect 10139 7644 10203 7648
rect 10139 7588 10143 7644
rect 10143 7588 10199 7644
rect 10199 7588 10203 7644
rect 10139 7584 10203 7588
rect 3114 7100 3178 7104
rect 3114 7044 3118 7100
rect 3118 7044 3174 7100
rect 3174 7044 3178 7100
rect 3114 7040 3178 7044
rect 3194 7100 3258 7104
rect 3194 7044 3198 7100
rect 3198 7044 3254 7100
rect 3254 7044 3258 7100
rect 3194 7040 3258 7044
rect 3274 7100 3338 7104
rect 3274 7044 3278 7100
rect 3278 7044 3334 7100
rect 3334 7044 3338 7100
rect 3274 7040 3338 7044
rect 3354 7100 3418 7104
rect 3354 7044 3358 7100
rect 3358 7044 3414 7100
rect 3414 7044 3418 7100
rect 3354 7040 3418 7044
rect 5828 7100 5892 7104
rect 5828 7044 5832 7100
rect 5832 7044 5888 7100
rect 5888 7044 5892 7100
rect 5828 7040 5892 7044
rect 5908 7100 5972 7104
rect 5908 7044 5912 7100
rect 5912 7044 5968 7100
rect 5968 7044 5972 7100
rect 5908 7040 5972 7044
rect 5988 7100 6052 7104
rect 5988 7044 5992 7100
rect 5992 7044 6048 7100
rect 6048 7044 6052 7100
rect 5988 7040 6052 7044
rect 6068 7100 6132 7104
rect 6068 7044 6072 7100
rect 6072 7044 6128 7100
rect 6128 7044 6132 7100
rect 6068 7040 6132 7044
rect 8542 7100 8606 7104
rect 8542 7044 8546 7100
rect 8546 7044 8602 7100
rect 8602 7044 8606 7100
rect 8542 7040 8606 7044
rect 8622 7100 8686 7104
rect 8622 7044 8626 7100
rect 8626 7044 8682 7100
rect 8682 7044 8686 7100
rect 8622 7040 8686 7044
rect 8702 7100 8766 7104
rect 8702 7044 8706 7100
rect 8706 7044 8762 7100
rect 8762 7044 8766 7100
rect 8702 7040 8766 7044
rect 8782 7100 8846 7104
rect 8782 7044 8786 7100
rect 8786 7044 8842 7100
rect 8842 7044 8846 7100
rect 8782 7040 8846 7044
rect 11256 7100 11320 7104
rect 11256 7044 11260 7100
rect 11260 7044 11316 7100
rect 11316 7044 11320 7100
rect 11256 7040 11320 7044
rect 11336 7100 11400 7104
rect 11336 7044 11340 7100
rect 11340 7044 11396 7100
rect 11396 7044 11400 7100
rect 11336 7040 11400 7044
rect 11416 7100 11480 7104
rect 11416 7044 11420 7100
rect 11420 7044 11476 7100
rect 11476 7044 11480 7100
rect 11416 7040 11480 7044
rect 11496 7100 11560 7104
rect 11496 7044 11500 7100
rect 11500 7044 11556 7100
rect 11556 7044 11560 7100
rect 11496 7040 11560 7044
rect 1757 6556 1821 6560
rect 1757 6500 1761 6556
rect 1761 6500 1817 6556
rect 1817 6500 1821 6556
rect 1757 6496 1821 6500
rect 1837 6556 1901 6560
rect 1837 6500 1841 6556
rect 1841 6500 1897 6556
rect 1897 6500 1901 6556
rect 1837 6496 1901 6500
rect 1917 6556 1981 6560
rect 1917 6500 1921 6556
rect 1921 6500 1977 6556
rect 1977 6500 1981 6556
rect 1917 6496 1981 6500
rect 1997 6556 2061 6560
rect 1997 6500 2001 6556
rect 2001 6500 2057 6556
rect 2057 6500 2061 6556
rect 1997 6496 2061 6500
rect 4471 6556 4535 6560
rect 4471 6500 4475 6556
rect 4475 6500 4531 6556
rect 4531 6500 4535 6556
rect 4471 6496 4535 6500
rect 4551 6556 4615 6560
rect 4551 6500 4555 6556
rect 4555 6500 4611 6556
rect 4611 6500 4615 6556
rect 4551 6496 4615 6500
rect 4631 6556 4695 6560
rect 4631 6500 4635 6556
rect 4635 6500 4691 6556
rect 4691 6500 4695 6556
rect 4631 6496 4695 6500
rect 4711 6556 4775 6560
rect 4711 6500 4715 6556
rect 4715 6500 4771 6556
rect 4771 6500 4775 6556
rect 4711 6496 4775 6500
rect 7185 6556 7249 6560
rect 7185 6500 7189 6556
rect 7189 6500 7245 6556
rect 7245 6500 7249 6556
rect 7185 6496 7249 6500
rect 7265 6556 7329 6560
rect 7265 6500 7269 6556
rect 7269 6500 7325 6556
rect 7325 6500 7329 6556
rect 7265 6496 7329 6500
rect 7345 6556 7409 6560
rect 7345 6500 7349 6556
rect 7349 6500 7405 6556
rect 7405 6500 7409 6556
rect 7345 6496 7409 6500
rect 7425 6556 7489 6560
rect 7425 6500 7429 6556
rect 7429 6500 7485 6556
rect 7485 6500 7489 6556
rect 7425 6496 7489 6500
rect 9899 6556 9963 6560
rect 9899 6500 9903 6556
rect 9903 6500 9959 6556
rect 9959 6500 9963 6556
rect 9899 6496 9963 6500
rect 9979 6556 10043 6560
rect 9979 6500 9983 6556
rect 9983 6500 10039 6556
rect 10039 6500 10043 6556
rect 9979 6496 10043 6500
rect 10059 6556 10123 6560
rect 10059 6500 10063 6556
rect 10063 6500 10119 6556
rect 10119 6500 10123 6556
rect 10059 6496 10123 6500
rect 10139 6556 10203 6560
rect 10139 6500 10143 6556
rect 10143 6500 10199 6556
rect 10199 6500 10203 6556
rect 10139 6496 10203 6500
rect 9076 6292 9140 6356
rect 3114 6012 3178 6016
rect 3114 5956 3118 6012
rect 3118 5956 3174 6012
rect 3174 5956 3178 6012
rect 3114 5952 3178 5956
rect 3194 6012 3258 6016
rect 3194 5956 3198 6012
rect 3198 5956 3254 6012
rect 3254 5956 3258 6012
rect 3194 5952 3258 5956
rect 3274 6012 3338 6016
rect 3274 5956 3278 6012
rect 3278 5956 3334 6012
rect 3334 5956 3338 6012
rect 3274 5952 3338 5956
rect 3354 6012 3418 6016
rect 3354 5956 3358 6012
rect 3358 5956 3414 6012
rect 3414 5956 3418 6012
rect 3354 5952 3418 5956
rect 5828 6012 5892 6016
rect 5828 5956 5832 6012
rect 5832 5956 5888 6012
rect 5888 5956 5892 6012
rect 5828 5952 5892 5956
rect 5908 6012 5972 6016
rect 5908 5956 5912 6012
rect 5912 5956 5968 6012
rect 5968 5956 5972 6012
rect 5908 5952 5972 5956
rect 5988 6012 6052 6016
rect 5988 5956 5992 6012
rect 5992 5956 6048 6012
rect 6048 5956 6052 6012
rect 5988 5952 6052 5956
rect 6068 6012 6132 6016
rect 6068 5956 6072 6012
rect 6072 5956 6128 6012
rect 6128 5956 6132 6012
rect 6068 5952 6132 5956
rect 8542 6012 8606 6016
rect 8542 5956 8546 6012
rect 8546 5956 8602 6012
rect 8602 5956 8606 6012
rect 8542 5952 8606 5956
rect 8622 6012 8686 6016
rect 8622 5956 8626 6012
rect 8626 5956 8682 6012
rect 8682 5956 8686 6012
rect 8622 5952 8686 5956
rect 8702 6012 8766 6016
rect 8702 5956 8706 6012
rect 8706 5956 8762 6012
rect 8762 5956 8766 6012
rect 8702 5952 8766 5956
rect 8782 6012 8846 6016
rect 8782 5956 8786 6012
rect 8786 5956 8842 6012
rect 8842 5956 8846 6012
rect 8782 5952 8846 5956
rect 11256 6012 11320 6016
rect 11256 5956 11260 6012
rect 11260 5956 11316 6012
rect 11316 5956 11320 6012
rect 11256 5952 11320 5956
rect 11336 6012 11400 6016
rect 11336 5956 11340 6012
rect 11340 5956 11396 6012
rect 11396 5956 11400 6012
rect 11336 5952 11400 5956
rect 11416 6012 11480 6016
rect 11416 5956 11420 6012
rect 11420 5956 11476 6012
rect 11476 5956 11480 6012
rect 11416 5952 11480 5956
rect 11496 6012 11560 6016
rect 11496 5956 11500 6012
rect 11500 5956 11556 6012
rect 11556 5956 11560 6012
rect 11496 5952 11560 5956
rect 1757 5468 1821 5472
rect 1757 5412 1761 5468
rect 1761 5412 1817 5468
rect 1817 5412 1821 5468
rect 1757 5408 1821 5412
rect 1837 5468 1901 5472
rect 1837 5412 1841 5468
rect 1841 5412 1897 5468
rect 1897 5412 1901 5468
rect 1837 5408 1901 5412
rect 1917 5468 1981 5472
rect 1917 5412 1921 5468
rect 1921 5412 1977 5468
rect 1977 5412 1981 5468
rect 1917 5408 1981 5412
rect 1997 5468 2061 5472
rect 1997 5412 2001 5468
rect 2001 5412 2057 5468
rect 2057 5412 2061 5468
rect 1997 5408 2061 5412
rect 4471 5468 4535 5472
rect 4471 5412 4475 5468
rect 4475 5412 4531 5468
rect 4531 5412 4535 5468
rect 4471 5408 4535 5412
rect 4551 5468 4615 5472
rect 4551 5412 4555 5468
rect 4555 5412 4611 5468
rect 4611 5412 4615 5468
rect 4551 5408 4615 5412
rect 4631 5468 4695 5472
rect 4631 5412 4635 5468
rect 4635 5412 4691 5468
rect 4691 5412 4695 5468
rect 4631 5408 4695 5412
rect 4711 5468 4775 5472
rect 4711 5412 4715 5468
rect 4715 5412 4771 5468
rect 4771 5412 4775 5468
rect 4711 5408 4775 5412
rect 7185 5468 7249 5472
rect 7185 5412 7189 5468
rect 7189 5412 7245 5468
rect 7245 5412 7249 5468
rect 7185 5408 7249 5412
rect 7265 5468 7329 5472
rect 7265 5412 7269 5468
rect 7269 5412 7325 5468
rect 7325 5412 7329 5468
rect 7265 5408 7329 5412
rect 7345 5468 7409 5472
rect 7345 5412 7349 5468
rect 7349 5412 7405 5468
rect 7405 5412 7409 5468
rect 7345 5408 7409 5412
rect 7425 5468 7489 5472
rect 7425 5412 7429 5468
rect 7429 5412 7485 5468
rect 7485 5412 7489 5468
rect 7425 5408 7489 5412
rect 9899 5468 9963 5472
rect 9899 5412 9903 5468
rect 9903 5412 9959 5468
rect 9959 5412 9963 5468
rect 9899 5408 9963 5412
rect 9979 5468 10043 5472
rect 9979 5412 9983 5468
rect 9983 5412 10039 5468
rect 10039 5412 10043 5468
rect 9979 5408 10043 5412
rect 10059 5468 10123 5472
rect 10059 5412 10063 5468
rect 10063 5412 10119 5468
rect 10119 5412 10123 5468
rect 10059 5408 10123 5412
rect 10139 5468 10203 5472
rect 10139 5412 10143 5468
rect 10143 5412 10199 5468
rect 10199 5412 10203 5468
rect 10139 5408 10203 5412
rect 3114 4924 3178 4928
rect 3114 4868 3118 4924
rect 3118 4868 3174 4924
rect 3174 4868 3178 4924
rect 3114 4864 3178 4868
rect 3194 4924 3258 4928
rect 3194 4868 3198 4924
rect 3198 4868 3254 4924
rect 3254 4868 3258 4924
rect 3194 4864 3258 4868
rect 3274 4924 3338 4928
rect 3274 4868 3278 4924
rect 3278 4868 3334 4924
rect 3334 4868 3338 4924
rect 3274 4864 3338 4868
rect 3354 4924 3418 4928
rect 3354 4868 3358 4924
rect 3358 4868 3414 4924
rect 3414 4868 3418 4924
rect 3354 4864 3418 4868
rect 5828 4924 5892 4928
rect 5828 4868 5832 4924
rect 5832 4868 5888 4924
rect 5888 4868 5892 4924
rect 5828 4864 5892 4868
rect 5908 4924 5972 4928
rect 5908 4868 5912 4924
rect 5912 4868 5968 4924
rect 5968 4868 5972 4924
rect 5908 4864 5972 4868
rect 5988 4924 6052 4928
rect 5988 4868 5992 4924
rect 5992 4868 6048 4924
rect 6048 4868 6052 4924
rect 5988 4864 6052 4868
rect 6068 4924 6132 4928
rect 6068 4868 6072 4924
rect 6072 4868 6128 4924
rect 6128 4868 6132 4924
rect 6068 4864 6132 4868
rect 8542 4924 8606 4928
rect 8542 4868 8546 4924
rect 8546 4868 8602 4924
rect 8602 4868 8606 4924
rect 8542 4864 8606 4868
rect 8622 4924 8686 4928
rect 8622 4868 8626 4924
rect 8626 4868 8682 4924
rect 8682 4868 8686 4924
rect 8622 4864 8686 4868
rect 8702 4924 8766 4928
rect 8702 4868 8706 4924
rect 8706 4868 8762 4924
rect 8762 4868 8766 4924
rect 8702 4864 8766 4868
rect 8782 4924 8846 4928
rect 8782 4868 8786 4924
rect 8786 4868 8842 4924
rect 8842 4868 8846 4924
rect 8782 4864 8846 4868
rect 11256 4924 11320 4928
rect 11256 4868 11260 4924
rect 11260 4868 11316 4924
rect 11316 4868 11320 4924
rect 11256 4864 11320 4868
rect 11336 4924 11400 4928
rect 11336 4868 11340 4924
rect 11340 4868 11396 4924
rect 11396 4868 11400 4924
rect 11336 4864 11400 4868
rect 11416 4924 11480 4928
rect 11416 4868 11420 4924
rect 11420 4868 11476 4924
rect 11476 4868 11480 4924
rect 11416 4864 11480 4868
rect 11496 4924 11560 4928
rect 11496 4868 11500 4924
rect 11500 4868 11556 4924
rect 11556 4868 11560 4924
rect 11496 4864 11560 4868
rect 1757 4380 1821 4384
rect 1757 4324 1761 4380
rect 1761 4324 1817 4380
rect 1817 4324 1821 4380
rect 1757 4320 1821 4324
rect 1837 4380 1901 4384
rect 1837 4324 1841 4380
rect 1841 4324 1897 4380
rect 1897 4324 1901 4380
rect 1837 4320 1901 4324
rect 1917 4380 1981 4384
rect 1917 4324 1921 4380
rect 1921 4324 1977 4380
rect 1977 4324 1981 4380
rect 1917 4320 1981 4324
rect 1997 4380 2061 4384
rect 1997 4324 2001 4380
rect 2001 4324 2057 4380
rect 2057 4324 2061 4380
rect 1997 4320 2061 4324
rect 4471 4380 4535 4384
rect 4471 4324 4475 4380
rect 4475 4324 4531 4380
rect 4531 4324 4535 4380
rect 4471 4320 4535 4324
rect 4551 4380 4615 4384
rect 4551 4324 4555 4380
rect 4555 4324 4611 4380
rect 4611 4324 4615 4380
rect 4551 4320 4615 4324
rect 4631 4380 4695 4384
rect 4631 4324 4635 4380
rect 4635 4324 4691 4380
rect 4691 4324 4695 4380
rect 4631 4320 4695 4324
rect 4711 4380 4775 4384
rect 4711 4324 4715 4380
rect 4715 4324 4771 4380
rect 4771 4324 4775 4380
rect 4711 4320 4775 4324
rect 7185 4380 7249 4384
rect 7185 4324 7189 4380
rect 7189 4324 7245 4380
rect 7245 4324 7249 4380
rect 7185 4320 7249 4324
rect 7265 4380 7329 4384
rect 7265 4324 7269 4380
rect 7269 4324 7325 4380
rect 7325 4324 7329 4380
rect 7265 4320 7329 4324
rect 7345 4380 7409 4384
rect 7345 4324 7349 4380
rect 7349 4324 7405 4380
rect 7405 4324 7409 4380
rect 7345 4320 7409 4324
rect 7425 4380 7489 4384
rect 7425 4324 7429 4380
rect 7429 4324 7485 4380
rect 7485 4324 7489 4380
rect 7425 4320 7489 4324
rect 9899 4380 9963 4384
rect 9899 4324 9903 4380
rect 9903 4324 9959 4380
rect 9959 4324 9963 4380
rect 9899 4320 9963 4324
rect 9979 4380 10043 4384
rect 9979 4324 9983 4380
rect 9983 4324 10039 4380
rect 10039 4324 10043 4380
rect 9979 4320 10043 4324
rect 10059 4380 10123 4384
rect 10059 4324 10063 4380
rect 10063 4324 10119 4380
rect 10119 4324 10123 4380
rect 10059 4320 10123 4324
rect 10139 4380 10203 4384
rect 10139 4324 10143 4380
rect 10143 4324 10199 4380
rect 10199 4324 10203 4380
rect 10139 4320 10203 4324
rect 3114 3836 3178 3840
rect 3114 3780 3118 3836
rect 3118 3780 3174 3836
rect 3174 3780 3178 3836
rect 3114 3776 3178 3780
rect 3194 3836 3258 3840
rect 3194 3780 3198 3836
rect 3198 3780 3254 3836
rect 3254 3780 3258 3836
rect 3194 3776 3258 3780
rect 3274 3836 3338 3840
rect 3274 3780 3278 3836
rect 3278 3780 3334 3836
rect 3334 3780 3338 3836
rect 3274 3776 3338 3780
rect 3354 3836 3418 3840
rect 3354 3780 3358 3836
rect 3358 3780 3414 3836
rect 3414 3780 3418 3836
rect 3354 3776 3418 3780
rect 5828 3836 5892 3840
rect 5828 3780 5832 3836
rect 5832 3780 5888 3836
rect 5888 3780 5892 3836
rect 5828 3776 5892 3780
rect 5908 3836 5972 3840
rect 5908 3780 5912 3836
rect 5912 3780 5968 3836
rect 5968 3780 5972 3836
rect 5908 3776 5972 3780
rect 5988 3836 6052 3840
rect 5988 3780 5992 3836
rect 5992 3780 6048 3836
rect 6048 3780 6052 3836
rect 5988 3776 6052 3780
rect 6068 3836 6132 3840
rect 6068 3780 6072 3836
rect 6072 3780 6128 3836
rect 6128 3780 6132 3836
rect 6068 3776 6132 3780
rect 8542 3836 8606 3840
rect 8542 3780 8546 3836
rect 8546 3780 8602 3836
rect 8602 3780 8606 3836
rect 8542 3776 8606 3780
rect 8622 3836 8686 3840
rect 8622 3780 8626 3836
rect 8626 3780 8682 3836
rect 8682 3780 8686 3836
rect 8622 3776 8686 3780
rect 8702 3836 8766 3840
rect 8702 3780 8706 3836
rect 8706 3780 8762 3836
rect 8762 3780 8766 3836
rect 8702 3776 8766 3780
rect 8782 3836 8846 3840
rect 8782 3780 8786 3836
rect 8786 3780 8842 3836
rect 8842 3780 8846 3836
rect 8782 3776 8846 3780
rect 11256 3836 11320 3840
rect 11256 3780 11260 3836
rect 11260 3780 11316 3836
rect 11316 3780 11320 3836
rect 11256 3776 11320 3780
rect 11336 3836 11400 3840
rect 11336 3780 11340 3836
rect 11340 3780 11396 3836
rect 11396 3780 11400 3836
rect 11336 3776 11400 3780
rect 11416 3836 11480 3840
rect 11416 3780 11420 3836
rect 11420 3780 11476 3836
rect 11476 3780 11480 3836
rect 11416 3776 11480 3780
rect 11496 3836 11560 3840
rect 11496 3780 11500 3836
rect 11500 3780 11556 3836
rect 11556 3780 11560 3836
rect 11496 3776 11560 3780
rect 1757 3292 1821 3296
rect 1757 3236 1761 3292
rect 1761 3236 1817 3292
rect 1817 3236 1821 3292
rect 1757 3232 1821 3236
rect 1837 3292 1901 3296
rect 1837 3236 1841 3292
rect 1841 3236 1897 3292
rect 1897 3236 1901 3292
rect 1837 3232 1901 3236
rect 1917 3292 1981 3296
rect 1917 3236 1921 3292
rect 1921 3236 1977 3292
rect 1977 3236 1981 3292
rect 1917 3232 1981 3236
rect 1997 3292 2061 3296
rect 1997 3236 2001 3292
rect 2001 3236 2057 3292
rect 2057 3236 2061 3292
rect 1997 3232 2061 3236
rect 4471 3292 4535 3296
rect 4471 3236 4475 3292
rect 4475 3236 4531 3292
rect 4531 3236 4535 3292
rect 4471 3232 4535 3236
rect 4551 3292 4615 3296
rect 4551 3236 4555 3292
rect 4555 3236 4611 3292
rect 4611 3236 4615 3292
rect 4551 3232 4615 3236
rect 4631 3292 4695 3296
rect 4631 3236 4635 3292
rect 4635 3236 4691 3292
rect 4691 3236 4695 3292
rect 4631 3232 4695 3236
rect 4711 3292 4775 3296
rect 4711 3236 4715 3292
rect 4715 3236 4771 3292
rect 4771 3236 4775 3292
rect 4711 3232 4775 3236
rect 7185 3292 7249 3296
rect 7185 3236 7189 3292
rect 7189 3236 7245 3292
rect 7245 3236 7249 3292
rect 7185 3232 7249 3236
rect 7265 3292 7329 3296
rect 7265 3236 7269 3292
rect 7269 3236 7325 3292
rect 7325 3236 7329 3292
rect 7265 3232 7329 3236
rect 7345 3292 7409 3296
rect 7345 3236 7349 3292
rect 7349 3236 7405 3292
rect 7405 3236 7409 3292
rect 7345 3232 7409 3236
rect 7425 3292 7489 3296
rect 7425 3236 7429 3292
rect 7429 3236 7485 3292
rect 7485 3236 7489 3292
rect 7425 3232 7489 3236
rect 9899 3292 9963 3296
rect 9899 3236 9903 3292
rect 9903 3236 9959 3292
rect 9959 3236 9963 3292
rect 9899 3232 9963 3236
rect 9979 3292 10043 3296
rect 9979 3236 9983 3292
rect 9983 3236 10039 3292
rect 10039 3236 10043 3292
rect 9979 3232 10043 3236
rect 10059 3292 10123 3296
rect 10059 3236 10063 3292
rect 10063 3236 10119 3292
rect 10119 3236 10123 3292
rect 10059 3232 10123 3236
rect 10139 3292 10203 3296
rect 10139 3236 10143 3292
rect 10143 3236 10199 3292
rect 10199 3236 10203 3292
rect 10139 3232 10203 3236
rect 3114 2748 3178 2752
rect 3114 2692 3118 2748
rect 3118 2692 3174 2748
rect 3174 2692 3178 2748
rect 3114 2688 3178 2692
rect 3194 2748 3258 2752
rect 3194 2692 3198 2748
rect 3198 2692 3254 2748
rect 3254 2692 3258 2748
rect 3194 2688 3258 2692
rect 3274 2748 3338 2752
rect 3274 2692 3278 2748
rect 3278 2692 3334 2748
rect 3334 2692 3338 2748
rect 3274 2688 3338 2692
rect 3354 2748 3418 2752
rect 3354 2692 3358 2748
rect 3358 2692 3414 2748
rect 3414 2692 3418 2748
rect 3354 2688 3418 2692
rect 5828 2748 5892 2752
rect 5828 2692 5832 2748
rect 5832 2692 5888 2748
rect 5888 2692 5892 2748
rect 5828 2688 5892 2692
rect 5908 2748 5972 2752
rect 5908 2692 5912 2748
rect 5912 2692 5968 2748
rect 5968 2692 5972 2748
rect 5908 2688 5972 2692
rect 5988 2748 6052 2752
rect 5988 2692 5992 2748
rect 5992 2692 6048 2748
rect 6048 2692 6052 2748
rect 5988 2688 6052 2692
rect 6068 2748 6132 2752
rect 6068 2692 6072 2748
rect 6072 2692 6128 2748
rect 6128 2692 6132 2748
rect 6068 2688 6132 2692
rect 8542 2748 8606 2752
rect 8542 2692 8546 2748
rect 8546 2692 8602 2748
rect 8602 2692 8606 2748
rect 8542 2688 8606 2692
rect 8622 2748 8686 2752
rect 8622 2692 8626 2748
rect 8626 2692 8682 2748
rect 8682 2692 8686 2748
rect 8622 2688 8686 2692
rect 8702 2748 8766 2752
rect 8702 2692 8706 2748
rect 8706 2692 8762 2748
rect 8762 2692 8766 2748
rect 8702 2688 8766 2692
rect 8782 2748 8846 2752
rect 8782 2692 8786 2748
rect 8786 2692 8842 2748
rect 8842 2692 8846 2748
rect 8782 2688 8846 2692
rect 11256 2748 11320 2752
rect 11256 2692 11260 2748
rect 11260 2692 11316 2748
rect 11316 2692 11320 2748
rect 11256 2688 11320 2692
rect 11336 2748 11400 2752
rect 11336 2692 11340 2748
rect 11340 2692 11396 2748
rect 11396 2692 11400 2748
rect 11336 2688 11400 2692
rect 11416 2748 11480 2752
rect 11416 2692 11420 2748
rect 11420 2692 11476 2748
rect 11476 2692 11480 2748
rect 11416 2688 11480 2692
rect 11496 2748 11560 2752
rect 11496 2692 11500 2748
rect 11500 2692 11556 2748
rect 11556 2692 11560 2748
rect 11496 2688 11560 2692
rect 1757 2204 1821 2208
rect 1757 2148 1761 2204
rect 1761 2148 1817 2204
rect 1817 2148 1821 2204
rect 1757 2144 1821 2148
rect 1837 2204 1901 2208
rect 1837 2148 1841 2204
rect 1841 2148 1897 2204
rect 1897 2148 1901 2204
rect 1837 2144 1901 2148
rect 1917 2204 1981 2208
rect 1917 2148 1921 2204
rect 1921 2148 1977 2204
rect 1977 2148 1981 2204
rect 1917 2144 1981 2148
rect 1997 2204 2061 2208
rect 1997 2148 2001 2204
rect 2001 2148 2057 2204
rect 2057 2148 2061 2204
rect 1997 2144 2061 2148
rect 4471 2204 4535 2208
rect 4471 2148 4475 2204
rect 4475 2148 4531 2204
rect 4531 2148 4535 2204
rect 4471 2144 4535 2148
rect 4551 2204 4615 2208
rect 4551 2148 4555 2204
rect 4555 2148 4611 2204
rect 4611 2148 4615 2204
rect 4551 2144 4615 2148
rect 4631 2204 4695 2208
rect 4631 2148 4635 2204
rect 4635 2148 4691 2204
rect 4691 2148 4695 2204
rect 4631 2144 4695 2148
rect 4711 2204 4775 2208
rect 4711 2148 4715 2204
rect 4715 2148 4771 2204
rect 4771 2148 4775 2204
rect 4711 2144 4775 2148
rect 7185 2204 7249 2208
rect 7185 2148 7189 2204
rect 7189 2148 7245 2204
rect 7245 2148 7249 2204
rect 7185 2144 7249 2148
rect 7265 2204 7329 2208
rect 7265 2148 7269 2204
rect 7269 2148 7325 2204
rect 7325 2148 7329 2204
rect 7265 2144 7329 2148
rect 7345 2204 7409 2208
rect 7345 2148 7349 2204
rect 7349 2148 7405 2204
rect 7405 2148 7409 2204
rect 7345 2144 7409 2148
rect 7425 2204 7489 2208
rect 7425 2148 7429 2204
rect 7429 2148 7485 2204
rect 7485 2148 7489 2204
rect 7425 2144 7489 2148
rect 9899 2204 9963 2208
rect 9899 2148 9903 2204
rect 9903 2148 9959 2204
rect 9959 2148 9963 2204
rect 9899 2144 9963 2148
rect 9979 2204 10043 2208
rect 9979 2148 9983 2204
rect 9983 2148 10039 2204
rect 10039 2148 10043 2204
rect 9979 2144 10043 2148
rect 10059 2204 10123 2208
rect 10059 2148 10063 2204
rect 10063 2148 10119 2204
rect 10119 2148 10123 2204
rect 10059 2144 10123 2148
rect 10139 2204 10203 2208
rect 10139 2148 10143 2204
rect 10143 2148 10199 2204
rect 10199 2148 10203 2204
rect 10139 2144 10203 2148
rect 3114 1660 3178 1664
rect 3114 1604 3118 1660
rect 3118 1604 3174 1660
rect 3174 1604 3178 1660
rect 3114 1600 3178 1604
rect 3194 1660 3258 1664
rect 3194 1604 3198 1660
rect 3198 1604 3254 1660
rect 3254 1604 3258 1660
rect 3194 1600 3258 1604
rect 3274 1660 3338 1664
rect 3274 1604 3278 1660
rect 3278 1604 3334 1660
rect 3334 1604 3338 1660
rect 3274 1600 3338 1604
rect 3354 1660 3418 1664
rect 3354 1604 3358 1660
rect 3358 1604 3414 1660
rect 3414 1604 3418 1660
rect 3354 1600 3418 1604
rect 5828 1660 5892 1664
rect 5828 1604 5832 1660
rect 5832 1604 5888 1660
rect 5888 1604 5892 1660
rect 5828 1600 5892 1604
rect 5908 1660 5972 1664
rect 5908 1604 5912 1660
rect 5912 1604 5968 1660
rect 5968 1604 5972 1660
rect 5908 1600 5972 1604
rect 5988 1660 6052 1664
rect 5988 1604 5992 1660
rect 5992 1604 6048 1660
rect 6048 1604 6052 1660
rect 5988 1600 6052 1604
rect 6068 1660 6132 1664
rect 6068 1604 6072 1660
rect 6072 1604 6128 1660
rect 6128 1604 6132 1660
rect 6068 1600 6132 1604
rect 8542 1660 8606 1664
rect 8542 1604 8546 1660
rect 8546 1604 8602 1660
rect 8602 1604 8606 1660
rect 8542 1600 8606 1604
rect 8622 1660 8686 1664
rect 8622 1604 8626 1660
rect 8626 1604 8682 1660
rect 8682 1604 8686 1660
rect 8622 1600 8686 1604
rect 8702 1660 8766 1664
rect 8702 1604 8706 1660
rect 8706 1604 8762 1660
rect 8762 1604 8766 1660
rect 8702 1600 8766 1604
rect 8782 1660 8846 1664
rect 8782 1604 8786 1660
rect 8786 1604 8842 1660
rect 8842 1604 8846 1660
rect 8782 1600 8846 1604
rect 11256 1660 11320 1664
rect 11256 1604 11260 1660
rect 11260 1604 11316 1660
rect 11316 1604 11320 1660
rect 11256 1600 11320 1604
rect 11336 1660 11400 1664
rect 11336 1604 11340 1660
rect 11340 1604 11396 1660
rect 11396 1604 11400 1660
rect 11336 1600 11400 1604
rect 11416 1660 11480 1664
rect 11416 1604 11420 1660
rect 11420 1604 11476 1660
rect 11476 1604 11480 1660
rect 11416 1600 11480 1604
rect 11496 1660 11560 1664
rect 11496 1604 11500 1660
rect 11500 1604 11556 1660
rect 11556 1604 11560 1660
rect 11496 1600 11560 1604
rect 1757 1116 1821 1120
rect 1757 1060 1761 1116
rect 1761 1060 1817 1116
rect 1817 1060 1821 1116
rect 1757 1056 1821 1060
rect 1837 1116 1901 1120
rect 1837 1060 1841 1116
rect 1841 1060 1897 1116
rect 1897 1060 1901 1116
rect 1837 1056 1901 1060
rect 1917 1116 1981 1120
rect 1917 1060 1921 1116
rect 1921 1060 1977 1116
rect 1977 1060 1981 1116
rect 1917 1056 1981 1060
rect 1997 1116 2061 1120
rect 1997 1060 2001 1116
rect 2001 1060 2057 1116
rect 2057 1060 2061 1116
rect 1997 1056 2061 1060
rect 4471 1116 4535 1120
rect 4471 1060 4475 1116
rect 4475 1060 4531 1116
rect 4531 1060 4535 1116
rect 4471 1056 4535 1060
rect 4551 1116 4615 1120
rect 4551 1060 4555 1116
rect 4555 1060 4611 1116
rect 4611 1060 4615 1116
rect 4551 1056 4615 1060
rect 4631 1116 4695 1120
rect 4631 1060 4635 1116
rect 4635 1060 4691 1116
rect 4691 1060 4695 1116
rect 4631 1056 4695 1060
rect 4711 1116 4775 1120
rect 4711 1060 4715 1116
rect 4715 1060 4771 1116
rect 4771 1060 4775 1116
rect 4711 1056 4775 1060
rect 7185 1116 7249 1120
rect 7185 1060 7189 1116
rect 7189 1060 7245 1116
rect 7245 1060 7249 1116
rect 7185 1056 7249 1060
rect 7265 1116 7329 1120
rect 7265 1060 7269 1116
rect 7269 1060 7325 1116
rect 7325 1060 7329 1116
rect 7265 1056 7329 1060
rect 7345 1116 7409 1120
rect 7345 1060 7349 1116
rect 7349 1060 7405 1116
rect 7405 1060 7409 1116
rect 7345 1056 7409 1060
rect 7425 1116 7489 1120
rect 7425 1060 7429 1116
rect 7429 1060 7485 1116
rect 7485 1060 7489 1116
rect 7425 1056 7489 1060
rect 9899 1116 9963 1120
rect 9899 1060 9903 1116
rect 9903 1060 9959 1116
rect 9959 1060 9963 1116
rect 9899 1056 9963 1060
rect 9979 1116 10043 1120
rect 9979 1060 9983 1116
rect 9983 1060 10039 1116
rect 10039 1060 10043 1116
rect 9979 1056 10043 1060
rect 10059 1116 10123 1120
rect 10059 1060 10063 1116
rect 10063 1060 10119 1116
rect 10119 1060 10123 1116
rect 10059 1056 10123 1060
rect 10139 1116 10203 1120
rect 10139 1060 10143 1116
rect 10143 1060 10199 1116
rect 10199 1060 10203 1116
rect 10139 1056 10203 1060
rect 3114 572 3178 576
rect 3114 516 3118 572
rect 3118 516 3174 572
rect 3174 516 3178 572
rect 3114 512 3178 516
rect 3194 572 3258 576
rect 3194 516 3198 572
rect 3198 516 3254 572
rect 3254 516 3258 572
rect 3194 512 3258 516
rect 3274 572 3338 576
rect 3274 516 3278 572
rect 3278 516 3334 572
rect 3334 516 3338 572
rect 3274 512 3338 516
rect 3354 572 3418 576
rect 3354 516 3358 572
rect 3358 516 3414 572
rect 3414 516 3418 572
rect 3354 512 3418 516
rect 5828 572 5892 576
rect 5828 516 5832 572
rect 5832 516 5888 572
rect 5888 516 5892 572
rect 5828 512 5892 516
rect 5908 572 5972 576
rect 5908 516 5912 572
rect 5912 516 5968 572
rect 5968 516 5972 572
rect 5908 512 5972 516
rect 5988 572 6052 576
rect 5988 516 5992 572
rect 5992 516 6048 572
rect 6048 516 6052 572
rect 5988 512 6052 516
rect 6068 572 6132 576
rect 6068 516 6072 572
rect 6072 516 6128 572
rect 6128 516 6132 572
rect 6068 512 6132 516
rect 8542 572 8606 576
rect 8542 516 8546 572
rect 8546 516 8602 572
rect 8602 516 8606 572
rect 8542 512 8606 516
rect 8622 572 8686 576
rect 8622 516 8626 572
rect 8626 516 8682 572
rect 8682 516 8686 572
rect 8622 512 8686 516
rect 8702 572 8766 576
rect 8702 516 8706 572
rect 8706 516 8762 572
rect 8762 516 8766 572
rect 8702 512 8766 516
rect 8782 572 8846 576
rect 8782 516 8786 572
rect 8786 516 8842 572
rect 8842 516 8846 572
rect 8782 512 8846 516
rect 11256 572 11320 576
rect 11256 516 11260 572
rect 11260 516 11316 572
rect 11316 516 11320 572
rect 11256 512 11320 516
rect 11336 572 11400 576
rect 11336 516 11340 572
rect 11340 516 11396 572
rect 11396 516 11400 572
rect 11336 512 11400 516
rect 11416 572 11480 576
rect 11416 516 11420 572
rect 11420 516 11476 572
rect 11476 516 11480 572
rect 11416 512 11480 516
rect 11496 572 11560 576
rect 11496 516 11500 572
rect 11500 516 11556 572
rect 11556 516 11560 572
rect 11496 512 11560 516
<< metal4 >>
rect 1749 10912 2069 11472
rect 1749 10848 1757 10912
rect 1821 10848 1837 10912
rect 1901 10848 1917 10912
rect 1981 10848 1997 10912
rect 2061 10848 2069 10912
rect 1749 9824 2069 10848
rect 1749 9760 1757 9824
rect 1821 9760 1837 9824
rect 1901 9760 1917 9824
rect 1981 9760 1997 9824
rect 2061 9760 2069 9824
rect 1749 8736 2069 9760
rect 1749 8672 1757 8736
rect 1821 8672 1837 8736
rect 1901 8672 1917 8736
rect 1981 8672 1997 8736
rect 2061 8672 2069 8736
rect 1749 7648 2069 8672
rect 1749 7584 1757 7648
rect 1821 7584 1837 7648
rect 1901 7584 1917 7648
rect 1981 7584 1997 7648
rect 2061 7584 2069 7648
rect 1749 6560 2069 7584
rect 1749 6496 1757 6560
rect 1821 6496 1837 6560
rect 1901 6496 1917 6560
rect 1981 6496 1997 6560
rect 2061 6496 2069 6560
rect 1749 5472 2069 6496
rect 1749 5408 1757 5472
rect 1821 5408 1837 5472
rect 1901 5408 1917 5472
rect 1981 5408 1997 5472
rect 2061 5408 2069 5472
rect 1749 4384 2069 5408
rect 1749 4320 1757 4384
rect 1821 4320 1837 4384
rect 1901 4320 1917 4384
rect 1981 4320 1997 4384
rect 2061 4320 2069 4384
rect 1749 3296 2069 4320
rect 1749 3232 1757 3296
rect 1821 3232 1837 3296
rect 1901 3232 1917 3296
rect 1981 3232 1997 3296
rect 2061 3232 2069 3296
rect 1749 2208 2069 3232
rect 1749 2144 1757 2208
rect 1821 2144 1837 2208
rect 1901 2144 1917 2208
rect 1981 2144 1997 2208
rect 2061 2144 2069 2208
rect 1749 1120 2069 2144
rect 1749 1056 1757 1120
rect 1821 1056 1837 1120
rect 1901 1056 1917 1120
rect 1981 1056 1997 1120
rect 2061 1056 2069 1120
rect 1749 496 2069 1056
rect 3106 11456 3426 11472
rect 3106 11392 3114 11456
rect 3178 11392 3194 11456
rect 3258 11392 3274 11456
rect 3338 11392 3354 11456
rect 3418 11392 3426 11456
rect 3106 10368 3426 11392
rect 3106 10304 3114 10368
rect 3178 10304 3194 10368
rect 3258 10304 3274 10368
rect 3338 10304 3354 10368
rect 3418 10304 3426 10368
rect 3106 9280 3426 10304
rect 3106 9216 3114 9280
rect 3178 9216 3194 9280
rect 3258 9216 3274 9280
rect 3338 9216 3354 9280
rect 3418 9216 3426 9280
rect 3106 8192 3426 9216
rect 3106 8128 3114 8192
rect 3178 8128 3194 8192
rect 3258 8128 3274 8192
rect 3338 8128 3354 8192
rect 3418 8128 3426 8192
rect 3106 7104 3426 8128
rect 3106 7040 3114 7104
rect 3178 7040 3194 7104
rect 3258 7040 3274 7104
rect 3338 7040 3354 7104
rect 3418 7040 3426 7104
rect 3106 6016 3426 7040
rect 3106 5952 3114 6016
rect 3178 5952 3194 6016
rect 3258 5952 3274 6016
rect 3338 5952 3354 6016
rect 3418 5952 3426 6016
rect 3106 4928 3426 5952
rect 3106 4864 3114 4928
rect 3178 4864 3194 4928
rect 3258 4864 3274 4928
rect 3338 4864 3354 4928
rect 3418 4864 3426 4928
rect 3106 3840 3426 4864
rect 3106 3776 3114 3840
rect 3178 3776 3194 3840
rect 3258 3776 3274 3840
rect 3338 3776 3354 3840
rect 3418 3776 3426 3840
rect 3106 2752 3426 3776
rect 3106 2688 3114 2752
rect 3178 2688 3194 2752
rect 3258 2688 3274 2752
rect 3338 2688 3354 2752
rect 3418 2688 3426 2752
rect 3106 1664 3426 2688
rect 3106 1600 3114 1664
rect 3178 1600 3194 1664
rect 3258 1600 3274 1664
rect 3338 1600 3354 1664
rect 3418 1600 3426 1664
rect 3106 576 3426 1600
rect 3106 512 3114 576
rect 3178 512 3194 576
rect 3258 512 3274 576
rect 3338 512 3354 576
rect 3418 512 3426 576
rect 3106 496 3426 512
rect 4463 10912 4783 11472
rect 4463 10848 4471 10912
rect 4535 10848 4551 10912
rect 4615 10848 4631 10912
rect 4695 10848 4711 10912
rect 4775 10848 4783 10912
rect 4463 9824 4783 10848
rect 4463 9760 4471 9824
rect 4535 9760 4551 9824
rect 4615 9760 4631 9824
rect 4695 9760 4711 9824
rect 4775 9760 4783 9824
rect 4463 8736 4783 9760
rect 4463 8672 4471 8736
rect 4535 8672 4551 8736
rect 4615 8672 4631 8736
rect 4695 8672 4711 8736
rect 4775 8672 4783 8736
rect 4463 7648 4783 8672
rect 4463 7584 4471 7648
rect 4535 7584 4551 7648
rect 4615 7584 4631 7648
rect 4695 7584 4711 7648
rect 4775 7584 4783 7648
rect 4463 6560 4783 7584
rect 4463 6496 4471 6560
rect 4535 6496 4551 6560
rect 4615 6496 4631 6560
rect 4695 6496 4711 6560
rect 4775 6496 4783 6560
rect 4463 5472 4783 6496
rect 4463 5408 4471 5472
rect 4535 5408 4551 5472
rect 4615 5408 4631 5472
rect 4695 5408 4711 5472
rect 4775 5408 4783 5472
rect 4463 4384 4783 5408
rect 4463 4320 4471 4384
rect 4535 4320 4551 4384
rect 4615 4320 4631 4384
rect 4695 4320 4711 4384
rect 4775 4320 4783 4384
rect 4463 3296 4783 4320
rect 4463 3232 4471 3296
rect 4535 3232 4551 3296
rect 4615 3232 4631 3296
rect 4695 3232 4711 3296
rect 4775 3232 4783 3296
rect 4463 2208 4783 3232
rect 4463 2144 4471 2208
rect 4535 2144 4551 2208
rect 4615 2144 4631 2208
rect 4695 2144 4711 2208
rect 4775 2144 4783 2208
rect 4463 1120 4783 2144
rect 4463 1056 4471 1120
rect 4535 1056 4551 1120
rect 4615 1056 4631 1120
rect 4695 1056 4711 1120
rect 4775 1056 4783 1120
rect 4463 496 4783 1056
rect 5820 11456 6140 11472
rect 5820 11392 5828 11456
rect 5892 11392 5908 11456
rect 5972 11392 5988 11456
rect 6052 11392 6068 11456
rect 6132 11392 6140 11456
rect 5820 10368 6140 11392
rect 5820 10304 5828 10368
rect 5892 10304 5908 10368
rect 5972 10304 5988 10368
rect 6052 10304 6068 10368
rect 6132 10304 6140 10368
rect 5820 9280 6140 10304
rect 5820 9216 5828 9280
rect 5892 9216 5908 9280
rect 5972 9216 5988 9280
rect 6052 9216 6068 9280
rect 6132 9216 6140 9280
rect 5820 8192 6140 9216
rect 5820 8128 5828 8192
rect 5892 8128 5908 8192
rect 5972 8128 5988 8192
rect 6052 8128 6068 8192
rect 6132 8128 6140 8192
rect 5820 7104 6140 8128
rect 5820 7040 5828 7104
rect 5892 7040 5908 7104
rect 5972 7040 5988 7104
rect 6052 7040 6068 7104
rect 6132 7040 6140 7104
rect 5820 6016 6140 7040
rect 5820 5952 5828 6016
rect 5892 5952 5908 6016
rect 5972 5952 5988 6016
rect 6052 5952 6068 6016
rect 6132 5952 6140 6016
rect 5820 4928 6140 5952
rect 5820 4864 5828 4928
rect 5892 4864 5908 4928
rect 5972 4864 5988 4928
rect 6052 4864 6068 4928
rect 6132 4864 6140 4928
rect 5820 3840 6140 4864
rect 5820 3776 5828 3840
rect 5892 3776 5908 3840
rect 5972 3776 5988 3840
rect 6052 3776 6068 3840
rect 6132 3776 6140 3840
rect 5820 2752 6140 3776
rect 5820 2688 5828 2752
rect 5892 2688 5908 2752
rect 5972 2688 5988 2752
rect 6052 2688 6068 2752
rect 6132 2688 6140 2752
rect 5820 1664 6140 2688
rect 5820 1600 5828 1664
rect 5892 1600 5908 1664
rect 5972 1600 5988 1664
rect 6052 1600 6068 1664
rect 6132 1600 6140 1664
rect 5820 576 6140 1600
rect 5820 512 5828 576
rect 5892 512 5908 576
rect 5972 512 5988 576
rect 6052 512 6068 576
rect 6132 512 6140 576
rect 5820 496 6140 512
rect 7177 10912 7497 11472
rect 7177 10848 7185 10912
rect 7249 10848 7265 10912
rect 7329 10848 7345 10912
rect 7409 10848 7425 10912
rect 7489 10848 7497 10912
rect 7177 9824 7497 10848
rect 7177 9760 7185 9824
rect 7249 9760 7265 9824
rect 7329 9760 7345 9824
rect 7409 9760 7425 9824
rect 7489 9760 7497 9824
rect 7177 8736 7497 9760
rect 7177 8672 7185 8736
rect 7249 8672 7265 8736
rect 7329 8672 7345 8736
rect 7409 8672 7425 8736
rect 7489 8672 7497 8736
rect 7177 7648 7497 8672
rect 7177 7584 7185 7648
rect 7249 7584 7265 7648
rect 7329 7584 7345 7648
rect 7409 7584 7425 7648
rect 7489 7584 7497 7648
rect 7177 6560 7497 7584
rect 7177 6496 7185 6560
rect 7249 6496 7265 6560
rect 7329 6496 7345 6560
rect 7409 6496 7425 6560
rect 7489 6496 7497 6560
rect 7177 5472 7497 6496
rect 7177 5408 7185 5472
rect 7249 5408 7265 5472
rect 7329 5408 7345 5472
rect 7409 5408 7425 5472
rect 7489 5408 7497 5472
rect 7177 4384 7497 5408
rect 7177 4320 7185 4384
rect 7249 4320 7265 4384
rect 7329 4320 7345 4384
rect 7409 4320 7425 4384
rect 7489 4320 7497 4384
rect 7177 3296 7497 4320
rect 7177 3232 7185 3296
rect 7249 3232 7265 3296
rect 7329 3232 7345 3296
rect 7409 3232 7425 3296
rect 7489 3232 7497 3296
rect 7177 2208 7497 3232
rect 7177 2144 7185 2208
rect 7249 2144 7265 2208
rect 7329 2144 7345 2208
rect 7409 2144 7425 2208
rect 7489 2144 7497 2208
rect 7177 1120 7497 2144
rect 7177 1056 7185 1120
rect 7249 1056 7265 1120
rect 7329 1056 7345 1120
rect 7409 1056 7425 1120
rect 7489 1056 7497 1120
rect 7177 496 7497 1056
rect 8534 11456 8854 11472
rect 8534 11392 8542 11456
rect 8606 11392 8622 11456
rect 8686 11392 8702 11456
rect 8766 11392 8782 11456
rect 8846 11392 8854 11456
rect 8534 10368 8854 11392
rect 8534 10304 8542 10368
rect 8606 10304 8622 10368
rect 8686 10304 8702 10368
rect 8766 10304 8782 10368
rect 8846 10304 8854 10368
rect 8534 9280 8854 10304
rect 9891 10912 10211 11472
rect 9891 10848 9899 10912
rect 9963 10848 9979 10912
rect 10043 10848 10059 10912
rect 10123 10848 10139 10912
rect 10203 10848 10211 10912
rect 9891 9824 10211 10848
rect 9891 9760 9899 9824
rect 9963 9760 9979 9824
rect 10043 9760 10059 9824
rect 10123 9760 10139 9824
rect 10203 9760 10211 9824
rect 9075 9620 9141 9621
rect 9075 9556 9076 9620
rect 9140 9556 9141 9620
rect 9075 9555 9141 9556
rect 8534 9216 8542 9280
rect 8606 9216 8622 9280
rect 8686 9216 8702 9280
rect 8766 9216 8782 9280
rect 8846 9216 8854 9280
rect 8534 8192 8854 9216
rect 8534 8128 8542 8192
rect 8606 8128 8622 8192
rect 8686 8128 8702 8192
rect 8766 8128 8782 8192
rect 8846 8128 8854 8192
rect 8534 7104 8854 8128
rect 8534 7040 8542 7104
rect 8606 7040 8622 7104
rect 8686 7040 8702 7104
rect 8766 7040 8782 7104
rect 8846 7040 8854 7104
rect 8534 6016 8854 7040
rect 9078 6357 9138 9555
rect 9891 8736 10211 9760
rect 9891 8672 9899 8736
rect 9963 8672 9979 8736
rect 10043 8672 10059 8736
rect 10123 8672 10139 8736
rect 10203 8672 10211 8736
rect 9891 7648 10211 8672
rect 9891 7584 9899 7648
rect 9963 7584 9979 7648
rect 10043 7584 10059 7648
rect 10123 7584 10139 7648
rect 10203 7584 10211 7648
rect 9891 6560 10211 7584
rect 9891 6496 9899 6560
rect 9963 6496 9979 6560
rect 10043 6496 10059 6560
rect 10123 6496 10139 6560
rect 10203 6496 10211 6560
rect 9075 6356 9141 6357
rect 9075 6292 9076 6356
rect 9140 6292 9141 6356
rect 9075 6291 9141 6292
rect 8534 5952 8542 6016
rect 8606 5952 8622 6016
rect 8686 5952 8702 6016
rect 8766 5952 8782 6016
rect 8846 5952 8854 6016
rect 8534 4928 8854 5952
rect 8534 4864 8542 4928
rect 8606 4864 8622 4928
rect 8686 4864 8702 4928
rect 8766 4864 8782 4928
rect 8846 4864 8854 4928
rect 8534 3840 8854 4864
rect 8534 3776 8542 3840
rect 8606 3776 8622 3840
rect 8686 3776 8702 3840
rect 8766 3776 8782 3840
rect 8846 3776 8854 3840
rect 8534 2752 8854 3776
rect 8534 2688 8542 2752
rect 8606 2688 8622 2752
rect 8686 2688 8702 2752
rect 8766 2688 8782 2752
rect 8846 2688 8854 2752
rect 8534 1664 8854 2688
rect 8534 1600 8542 1664
rect 8606 1600 8622 1664
rect 8686 1600 8702 1664
rect 8766 1600 8782 1664
rect 8846 1600 8854 1664
rect 8534 576 8854 1600
rect 8534 512 8542 576
rect 8606 512 8622 576
rect 8686 512 8702 576
rect 8766 512 8782 576
rect 8846 512 8854 576
rect 8534 496 8854 512
rect 9891 5472 10211 6496
rect 9891 5408 9899 5472
rect 9963 5408 9979 5472
rect 10043 5408 10059 5472
rect 10123 5408 10139 5472
rect 10203 5408 10211 5472
rect 9891 4384 10211 5408
rect 9891 4320 9899 4384
rect 9963 4320 9979 4384
rect 10043 4320 10059 4384
rect 10123 4320 10139 4384
rect 10203 4320 10211 4384
rect 9891 3296 10211 4320
rect 9891 3232 9899 3296
rect 9963 3232 9979 3296
rect 10043 3232 10059 3296
rect 10123 3232 10139 3296
rect 10203 3232 10211 3296
rect 9891 2208 10211 3232
rect 9891 2144 9899 2208
rect 9963 2144 9979 2208
rect 10043 2144 10059 2208
rect 10123 2144 10139 2208
rect 10203 2144 10211 2208
rect 9891 1120 10211 2144
rect 9891 1056 9899 1120
rect 9963 1056 9979 1120
rect 10043 1056 10059 1120
rect 10123 1056 10139 1120
rect 10203 1056 10211 1120
rect 9891 496 10211 1056
rect 11248 11456 11568 11472
rect 11248 11392 11256 11456
rect 11320 11392 11336 11456
rect 11400 11392 11416 11456
rect 11480 11392 11496 11456
rect 11560 11392 11568 11456
rect 11248 10368 11568 11392
rect 11248 10304 11256 10368
rect 11320 10304 11336 10368
rect 11400 10304 11416 10368
rect 11480 10304 11496 10368
rect 11560 10304 11568 10368
rect 11248 9280 11568 10304
rect 11248 9216 11256 9280
rect 11320 9216 11336 9280
rect 11400 9216 11416 9280
rect 11480 9216 11496 9280
rect 11560 9216 11568 9280
rect 11248 8192 11568 9216
rect 11248 8128 11256 8192
rect 11320 8128 11336 8192
rect 11400 8128 11416 8192
rect 11480 8128 11496 8192
rect 11560 8128 11568 8192
rect 11248 7104 11568 8128
rect 11248 7040 11256 7104
rect 11320 7040 11336 7104
rect 11400 7040 11416 7104
rect 11480 7040 11496 7104
rect 11560 7040 11568 7104
rect 11248 6016 11568 7040
rect 11248 5952 11256 6016
rect 11320 5952 11336 6016
rect 11400 5952 11416 6016
rect 11480 5952 11496 6016
rect 11560 5952 11568 6016
rect 11248 4928 11568 5952
rect 11248 4864 11256 4928
rect 11320 4864 11336 4928
rect 11400 4864 11416 4928
rect 11480 4864 11496 4928
rect 11560 4864 11568 4928
rect 11248 3840 11568 4864
rect 11248 3776 11256 3840
rect 11320 3776 11336 3840
rect 11400 3776 11416 3840
rect 11480 3776 11496 3840
rect 11560 3776 11568 3840
rect 11248 2752 11568 3776
rect 11248 2688 11256 2752
rect 11320 2688 11336 2752
rect 11400 2688 11416 2752
rect 11480 2688 11496 2752
rect 11560 2688 11568 2752
rect 11248 1664 11568 2688
rect 11248 1600 11256 1664
rect 11320 1600 11336 1664
rect 11400 1600 11416 1664
rect 11480 1600 11496 1664
rect 11560 1600 11568 1664
rect 11248 576 11568 1600
rect 11248 512 11256 576
rect 11320 512 11336 576
rect 11400 512 11416 576
rect 11480 512 11496 576
rect 11560 512 11568 576
rect 11248 496 11568 512
use sky130_fd_sc_hd__and4_1  _065_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 4968 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _066_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 7268 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _067_
timestamp 1701704242
transform 1 0 8096 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _068_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 9292 0 1 7072
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _069_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 3128 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _070_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 9476 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _071_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 9660 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _072_
timestamp 1701704242
transform 1 0 10488 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _073_
timestamp 1701704242
transform -1 0 10856 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _074_
timestamp 1701704242
transform 1 0 9936 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _075_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 10856 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1701704242
transform -1 0 8924 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _077_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 10856 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _078_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 8924 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _079_
timestamp 1701704242
transform 1 0 8924 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _080_
timestamp 1701704242
transform -1 0 10856 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _081_
timestamp 1701704242
transform -1 0 10580 0 -1 10336
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _082_
timestamp 1701704242
transform 1 0 10580 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _083_
timestamp 1701704242
transform 1 0 8004 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _084_
timestamp 1701704242
transform 1 0 5244 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _085_
timestamp 1701704242
transform -1 0 8924 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _086_
timestamp 1701704242
transform -1 0 8280 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _087_
timestamp 1701704242
transform -1 0 8280 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _088_
timestamp 1701704242
transform -1 0 7912 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _089_
timestamp 1701704242
transform -1 0 7544 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _090_
timestamp 1701704242
transform 1 0 6716 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _091_
timestamp 1701704242
transform 1 0 7544 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _092_
timestamp 1701704242
transform 1 0 5796 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _093_
timestamp 1701704242
transform -1 0 7728 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _094_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 5980 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _095_
timestamp 1701704242
transform -1 0 5152 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _096_
timestamp 1701704242
transform 1 0 5152 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _097_
timestamp 1701704242
transform -1 0 4232 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _098_
timestamp 1701704242
transform 1 0 4968 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _099_
timestamp 1701704242
transform -1 0 3588 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _100_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3588 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _101_
timestamp 1701704242
transform -1 0 1288 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _102_
timestamp 1701704242
transform 1 0 3220 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _103_
timestamp 1701704242
transform -1 0 3680 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _104_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3128 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 2300 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _106_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 2852 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _107_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 1288 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _108_
timestamp 1701704242
transform 1 0 2392 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _109_
timestamp 1701704242
transform -1 0 1656 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _110_
timestamp 1701704242
transform -1 0 5244 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _111_
timestamp 1701704242
transform -1 0 3496 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _112_
timestamp 1701704242
transform 1 0 3680 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _113_
timestamp 1701704242
transform 1 0 2576 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _114_
timestamp 1701704242
transform 1 0 3220 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _115_
timestamp 1701704242
transform -1 0 5520 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _116_
timestamp 1701704242
transform -1 0 3864 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _117_
timestamp 1701704242
transform -1 0 5428 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _118_
timestamp 1701704242
transform 1 0 4140 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _119_
timestamp 1701704242
transform 1 0 7084 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _120_
timestamp 1701704242
transform -1 0 6348 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _121_
timestamp 1701704242
transform 1 0 5980 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _122_
timestamp 1701704242
transform -1 0 7452 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _123_
timestamp 1701704242
transform 1 0 7728 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _124_
timestamp 1701704242
transform -1 0 8188 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _125_
timestamp 1701704242
transform 1 0 7452 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _126_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 6532 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _127_
timestamp 1701704242
transform 1 0 9292 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _128_
timestamp 1701704242
transform 1 0 8372 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _129_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 9292 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _130_
timestamp 1701704242
transform -1 0 10948 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _131_
timestamp 1701704242
transform 1 0 8924 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _132_
timestamp 1701704242
transform 1 0 8924 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _133_
timestamp 1701704242
transform 1 0 8372 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _134_
timestamp 1701704242
transform 1 0 7084 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _135_
timestamp 1701704242
transform 1 0 5612 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _136_
timestamp 1701704242
transform 1 0 5244 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _137_
timestamp 1701704242
transform -1 0 4876 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _138_
timestamp 1701704242
transform 1 0 3404 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _139_
timestamp 1701704242
transform -1 0 3128 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _140_
timestamp 1701704242
transform -1 0 2760 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _141__2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 10856 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _141_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 11132 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _142_
timestamp 1701704242
transform 1 0 3128 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _143_
timestamp 1701704242
transform 1 0 2208 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _144_
timestamp 1701704242
transform 1 0 3680 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _145_
timestamp 1701704242
transform 1 0 3680 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _146_
timestamp 1701704242
transform 1 0 5612 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _147_
timestamp 1701704242
transform 1 0 5796 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _148_
timestamp 1701704242
transform 1 0 6348 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _149_
timestamp 1701704242
transform 1 0 7820 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _151_
timestamp 1701704242
transform -1 0 5244 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _152_
timestamp 1701704242
transform -1 0 6716 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _153_
timestamp 1701704242
transform 1 0 9292 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _154_
timestamp 1701704242
transform -1 0 6348 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _155_
timestamp 1701704242
transform 1 0 3864 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _156_
timestamp 1701704242
transform -1 0 3128 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _157_
timestamp 1701704242
transform -1 0 1932 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _158_
timestamp 1701704242
transform -1 0 1564 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 7912 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1701704242
transform -1 0 5520 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1701704242
transform 1 0 8556 0 -1 9248
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1701704242
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1701704242
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1701704242
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1701704242
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1701704242
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1701704242
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1701704242
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1701704242
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1701704242
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10948 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1701704242
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1701704242
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1701704242
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1701704242
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1701704242
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1701704242
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1701704242
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1701704242
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1701704242
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1701704242
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_113
timestamp 1701704242
transform 1 0 10948 0 -1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1701704242
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1701704242
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1701704242
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1701704242
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1701704242
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1701704242
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1701704242
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1701704242
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1701704242
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1701704242
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1701704242
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_109
timestamp 1701704242
transform 1 0 10580 0 1 1632
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1701704242
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1701704242
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1701704242
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1701704242
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1701704242
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1701704242
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1701704242
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1701704242
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1701704242
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1701704242
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1701704242
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1701704242
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_113
timestamp 1701704242
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1701704242
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1701704242
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1701704242
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1701704242
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1701704242
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1701704242
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1701704242
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1701704242
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1701704242
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1701704242
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1701704242
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_109
timestamp 1701704242
transform 1 0 10580 0 1 2720
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1701704242
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1701704242
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1701704242
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1701704242
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1701704242
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1701704242
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1701704242
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1701704242
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1701704242
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1701704242
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1701704242
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1701704242
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_113
timestamp 1701704242
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1701704242
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1701704242
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1701704242
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1701704242
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1701704242
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1701704242
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1701704242
transform 1 0 6532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1701704242
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1701704242
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1701704242
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1701704242
transform 1 0 9476 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_109
timestamp 1701704242
transform 1 0 10580 0 1 3808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1701704242
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1701704242
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1701704242
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1701704242
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1701704242
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1701704242
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1701704242
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1701704242
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1701704242
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1701704242
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_105
timestamp 1701704242
transform 1 0 10212 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_113
timestamp 1701704242
transform 1 0 10948 0 -1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1701704242
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1701704242
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1701704242
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1701704242
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1701704242
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1701704242
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1701704242
transform 1 0 6532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1701704242
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1701704242
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1701704242
transform 1 0 8372 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_97
timestamp 1701704242
transform 1 0 9476 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_101
timestamp 1701704242
transform 1 0 9844 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_112
timestamp 1701704242
transform 1 0 10856 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1701704242
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1701704242
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1701704242
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1701704242
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1701704242
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1701704242
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1701704242
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_69
timestamp 1701704242
transform 1 0 6900 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_78 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 7728 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_86
timestamp 1701704242
transform 1 0 8464 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_91
timestamp 1701704242
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_97
timestamp 1701704242
transform 1 0 9476 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_113
timestamp 1701704242
transform 1 0 10948 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1701704242
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1701704242
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1701704242
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_29
timestamp 1701704242
transform 1 0 3220 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_33
timestamp 1701704242
transform 1 0 3588 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_38
timestamp 1701704242
transform 1 0 4048 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_45
timestamp 1701704242
transform 1 0 4692 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_55
timestamp 1701704242
transform 1 0 5612 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_73
timestamp 1701704242
transform 1 0 7268 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1701704242
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_85
timestamp 1701704242
transform 1 0 8372 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_113
timestamp 1701704242
transform 1 0 10948 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1701704242
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_15
timestamp 1701704242
transform 1 0 1932 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_53
timestamp 1701704242
transform 1 0 5428 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_57
timestamp 1701704242
transform 1 0 5796 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1701704242
transform 1 0 10764 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_113
timestamp 1701704242
transform 1 0 10948 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_3
timestamp 1701704242
transform 1 0 828 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_11
timestamp 1701704242
transform 1 0 1564 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_54
timestamp 1701704242
transform 1 0 5520 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_75
timestamp 1701704242
transform 1 0 7452 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_114
timestamp 1701704242
transform 1 0 11040 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1701704242
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_15
timestamp 1701704242
transform 1 0 1932 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_21
timestamp 1701704242
transform 1 0 2484 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_44
timestamp 1701704242
transform 1 0 4600 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_54
timestamp 1701704242
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_65
timestamp 1701704242
transform 1 0 6532 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_89
timestamp 1701704242
transform 1 0 8740 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_113
timestamp 1701704242
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1701704242
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_15
timestamp 1701704242
transform 1 0 1932 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_23
timestamp 1701704242
transform 1 0 2668 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_76
timestamp 1701704242
transform 1 0 7544 0 1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1701704242
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_15
timestamp 1701704242
transform 1 0 1932 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_19
timestamp 1701704242
transform 1 0 2300 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_27
timestamp 1701704242
transform 1 0 3036 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 1701704242
transform 1 0 5520 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_80
timestamp 1701704242
transform 1 0 7912 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_113
timestamp 1701704242
transform 1 0 10948 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_3
timestamp 1701704242
transform 1 0 828 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_29
timestamp 1701704242
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1701704242
transform 1 0 8188 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_3
timestamp 1701704242
transform 1 0 828 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_113
timestamp 1701704242
transform 1 0 10948 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_3
timestamp 1701704242
transform 1 0 828 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_23
timestamp 1701704242
transform 1 0 2668 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_93
timestamp 1701704242
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1701704242
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_15
timestamp 1701704242
transform 1 0 1932 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_26
timestamp 1701704242
transform 1 0 2944 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_54
timestamp 1701704242
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_57
timestamp 1701704242
transform 1 0 5796 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_113
timestamp 1701704242
transform 1 0 10948 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 5612 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1701704242
transform -1 0 9660 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1701704242
transform -1 0 11132 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1701704242
transform -1 0 11132 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1701704242
transform 1 0 1932 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1701704242
transform -1 0 7452 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1701704242
transform -1 0 4968 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1701704242
transform -1 0 7084 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1701704242
transform 1 0 9752 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1701704242
transform 1 0 10304 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1701704242
transform -1 0 6532 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1701704242
transform -1 0 5520 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1701704242
transform -1 0 9108 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1701704242
transform -1 0 9292 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1701704242
transform -1 0 10304 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1701704242
transform 1 0 7452 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1701704242
transform -1 0 3128 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1701704242
transform 1 0 1656 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1701704242
transform -1 0 7452 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1701704242
transform -1 0 10580 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1701704242
transform -1 0 4968 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1701704242
transform 1 0 4232 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1701704242
transform 1 0 7544 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1701704242
transform 1 0 5796 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_20
timestamp 1701704242
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1701704242
transform -1 0 11408 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_21
timestamp 1701704242
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1701704242
transform -1 0 11408 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_22
timestamp 1701704242
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1701704242
transform -1 0 11408 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_23
timestamp 1701704242
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1701704242
transform -1 0 11408 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_24
timestamp 1701704242
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1701704242
transform -1 0 11408 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_25
timestamp 1701704242
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1701704242
transform -1 0 11408 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_26
timestamp 1701704242
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1701704242
transform -1 0 11408 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_27
timestamp 1701704242
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1701704242
transform -1 0 11408 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_28
timestamp 1701704242
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1701704242
transform -1 0 11408 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_29
timestamp 1701704242
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1701704242
transform -1 0 11408 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_30
timestamp 1701704242
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1701704242
transform -1 0 11408 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_31
timestamp 1701704242
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1701704242
transform -1 0 11408 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_32
timestamp 1701704242
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1701704242
transform -1 0 11408 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_33
timestamp 1701704242
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1701704242
transform -1 0 11408 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_34
timestamp 1701704242
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1701704242
transform -1 0 11408 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_35
timestamp 1701704242
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1701704242
transform -1 0 11408 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_36
timestamp 1701704242
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1701704242
transform -1 0 11408 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_37
timestamp 1701704242
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1701704242
transform -1 0 11408 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_38
timestamp 1701704242
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1701704242
transform -1 0 11408 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_39
timestamp 1701704242
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1701704242
transform -1 0 11408 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_40 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_41
timestamp 1701704242
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_42
timestamp 1701704242
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_43
timestamp 1701704242
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_44
timestamp 1701704242
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_45
timestamp 1701704242
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_46
timestamp 1701704242
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_47
timestamp 1701704242
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_48
timestamp 1701704242
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_49
timestamp 1701704242
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_50
timestamp 1701704242
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_51
timestamp 1701704242
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_52
timestamp 1701704242
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_53
timestamp 1701704242
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_54
timestamp 1701704242
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_55
timestamp 1701704242
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_56
timestamp 1701704242
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_57
timestamp 1701704242
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_58
timestamp 1701704242
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_59
timestamp 1701704242
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_60
timestamp 1701704242
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_61
timestamp 1701704242
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_62
timestamp 1701704242
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_63
timestamp 1701704242
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_64
timestamp 1701704242
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_65
timestamp 1701704242
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_66
timestamp 1701704242
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_67
timestamp 1701704242
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_68
timestamp 1701704242
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_69
timestamp 1701704242
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_70
timestamp 1701704242
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_71
timestamp 1701704242
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_72
timestamp 1701704242
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_73
timestamp 1701704242
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_74
timestamp 1701704242
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_75
timestamp 1701704242
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_76
timestamp 1701704242
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_77
timestamp 1701704242
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_78
timestamp 1701704242
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_79
timestamp 1701704242
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_80
timestamp 1701704242
transform 1 0 3128 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_81
timestamp 1701704242
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_82
timestamp 1701704242
transform 1 0 8280 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_83
timestamp 1701704242
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
<< labels >>
rlabel metal2 s 6060 11424 6060 11424 4 VGND
rlabel metal1 s 5980 10880 5980 10880 4 VPWR
rlabel metal1 s 5842 10438 5842 10438 4 _000_
rlabel metal2 s 9609 6834 9609 6834 4 _001_
rlabel metal1 s 10733 6154 10733 6154 4 _002_
rlabel metal1 s 9016 6426 9016 6426 4 _003_
rlabel metal1 s 8556 9146 8556 9146 4 _004_
rlabel metal1 s 8924 9690 8924 9690 4 _005_
rlabel metal1 s 7539 10098 7539 10098 4 _006_
rlabel metal2 s 5842 9777 5842 9777 4 _007_
rlabel metal1 s 5290 10234 5290 10234 4 _008_
rlabel metal1 s 4799 10166 4799 10166 4 _009_
rlabel metal3 s 2300 9588 2300 9588 4 _010_
rlabel metal1 s 2852 8602 2852 8602 4 _011_
rlabel metal1 s 2028 9486 2028 9486 4 _012_
rlabel metal2 s 3445 7922 3445 7922 4 _013_
rlabel metal1 s 2208 7378 2208 7378 4 _014_
rlabel metal1 s 3900 7310 3900 7310 4 _015_
rlabel metal1 s 4094 6426 4094 6426 4 _016_
rlabel metal1 s 6067 7310 6067 7310 4 _017_
rlabel metal1 s 6481 6222 6481 6222 4 _018_
rlabel metal2 s 6665 6834 6665 6834 4 _019_
rlabel metal1 s 8275 6834 8275 6834 4 _020_
rlabel metal2 s 7958 7956 7958 7956 4 _021_
rlabel metal2 s 7774 8976 7774 8976 4 _022_
rlabel metal1 s 7222 8058 7222 8058 4 _023_
rlabel metal2 s 9338 7888 9338 7888 4 _024_
rlabel metal1 s 5658 8398 5658 8398 4 _025_
rlabel metal1 s 8096 7990 8096 7990 4 _026_
rlabel metal2 s 9246 7548 9246 7548 4 _027_
rlabel metal1 s 10304 7922 10304 7922 4 _028_
rlabel metal1 s 3680 9690 3680 9690 4 _029_
rlabel metal2 s 9430 6766 9430 6766 4 _030_
rlabel metal2 s 10534 6460 10534 6460 4 _031_
rlabel metal2 s 10442 8398 10442 8398 4 _032_
rlabel metal2 s 10350 5746 10350 5746 4 _033_
rlabel metal1 s 4140 10574 4140 10574 4 _034_
rlabel metal1 s 8878 5780 8878 5780 4 _035_
rlabel metal1 s 8970 5882 8970 5882 4 _036_
rlabel metal1 s 10396 8058 10396 8058 4 _037_
rlabel metal1 s 10258 9996 10258 9996 4 _038_
rlabel metal1 s 8234 8976 8234 8976 4 _039_
rlabel metal1 s 5934 9690 5934 9690 4 _040_
rlabel metal2 s 8234 10404 8234 10404 4 _041_
rlabel metal1 s 7728 10574 7728 10574 4 _042_
rlabel metal1 s 7314 10438 7314 10438 4 _043_
rlabel metal1 s 6348 11050 6348 11050 4 _044_
rlabel metal1 s 6440 10098 6440 10098 4 _045_
rlabel metal1 s 5842 8432 5842 8432 4 _046_
rlabel metal1 s 3404 10098 3404 10098 4 _047_
rlabel metal1 s 5382 10064 5382 10064 4 _048_
rlabel metal2 s 5198 9860 5198 9860 4 _049_
rlabel metal2 s 1058 10404 1058 10404 4 _050_
rlabel metal2 s 1242 10302 1242 10302 4 _051_
rlabel metal1 s 2714 11016 2714 11016 4 _052_
rlabel metal1 s 2691 9010 2691 9010 4 _053_
rlabel metal1 s 1518 10166 1518 10166 4 _054_
rlabel metal1 s 3036 8398 3036 8398 4 _055_
rlabel metal2 s 1150 9894 1150 9894 4 _056_
rlabel metal2 s 2438 9622 2438 9622 4 _057_
rlabel metal2 s 2806 7174 2806 7174 4 _058_
rlabel metal2 s 3634 6766 3634 6766 4 _059_
rlabel metal2 s 5474 7684 5474 7684 4 _060_
rlabel metal1 s 4370 6256 4370 6256 4 _061_
rlabel metal2 s 7130 7106 7130 7106 4 _062_
rlabel metal2 s 6302 7548 6302 7548 4 _063_
rlabel metal2 s 7866 7395 7866 7395 4 clk
rlabel metal1 s 6578 9112 6578 9112 4 clknet_0_clk
rlabel metal1 s 3496 9486 3496 9486 4 clknet_1_0__leaf_clk
rlabel metal1 s 10718 9078 10718 9078 4 clknet_1_1__leaf_clk
rlabel metal1 s 5244 9622 5244 9622 4 count[0]
rlabel metal1 s 7406 11322 7406 11322 4 count[1]
rlabel metal2 s 9522 10880 9522 10880 4 count[2]
rlabel metal1 s 6164 11322 6164 11322 4 count[3]
rlabel metal1 s 4370 11322 4370 11322 4 count[4]
rlabel metal2 s 2898 11152 2898 11152 4 count[5]
rlabel metal1 s 1932 10778 1932 10778 4 count[6]
rlabel metal1 s 1058 10778 1058 10778 4 count[7]
rlabel metal1 s 3128 7242 3128 7242 4 counter\[0\]
rlabel metal1 s 10902 7786 10902 7786 4 counter\[10\]
rlabel metal1 s 10994 9588 10994 9588 4 counter\[11\]
rlabel metal1 s 8004 10438 8004 10438 4 counter\[12\]
rlabel metal2 s 8050 11390 8050 11390 4 counter\[13\]
rlabel metal2 s 7038 10608 7038 10608 4 counter\[14\]
rlabel metal1 s 7452 10574 7452 10574 4 counter\[15\]
rlabel metal1 s 3818 9078 3818 9078 4 counter\[16\]
rlabel metal1 s 4462 9350 4462 9350 4 counter\[17\]
rlabel metal1 s 2300 10574 2300 10574 4 counter\[18\]
rlabel metal1 s 1426 10574 1426 10574 4 counter\[19\]
rlabel metal2 s 5198 7786 5198 7786 4 counter\[1\]
rlabel metal1 s 5106 7208 5106 7208 4 counter\[2\]
rlabel metal2 s 5106 7514 5106 7514 4 counter\[3\]
rlabel metal1 s 7866 7888 7866 7888 4 counter\[4\]
rlabel metal2 s 7590 7106 7590 7106 4 counter\[5\]
rlabel metal2 s 7774 6188 7774 6188 4 counter\[6\]
rlabel metal1 s 8924 7854 8924 7854 4 counter\[7\]
rlabel metal1 s 10764 6970 10764 6970 4 counter\[8\]
rlabel metal2 s 9890 6426 9890 6426 4 counter\[9\]
rlabel metal1 s 6210 9010 6210 9010 4 n_rst
rlabel metal1 s 5796 9146 5796 9146 4 net1
rlabel metal1 s 6348 10030 6348 10030 4 net10
rlabel metal1 s 10488 5746 10488 5746 4 net11
rlabel metal2 s 10718 5916 10718 5916 4 net12
rlabel metal1 s 5520 7310 5520 7310 4 net13
rlabel metal1 s 4784 8058 4784 8058 4 net14
rlabel metal1 s 8326 10506 8326 10506 4 net15
rlabel metal1 s 8372 10234 8372 10234 4 net16
rlabel metal1 s 9430 7174 9430 7174 4 net17
rlabel metal2 s 8142 7191 8142 7191 4 net18
rlabel metal2 s 2990 7616 2990 7616 4 net19
rlabel metal2 s 10810 10880 10810 10880 4 net2
rlabel metal2 s 2525 6834 2525 6834 4 net20
rlabel metal1 s 6624 8058 6624 8058 4 net21
rlabel metal1 s 8418 9418 8418 9418 4 net22
rlabel metal1 s 3910 10506 3910 10506 4 net23
rlabel metal1 s 5198 11118 5198 11118 4 net24
rlabel metal2 s 8234 7684 8234 7684 4 net25
rlabel metal1 s 4784 6222 4784 6222 4 net3
rlabel metal2 s 8970 8211 8970 8211 4 net4
rlabel metal1 s 9476 9010 9476 9010 4 net5
rlabel metal1 s 9476 6290 9476 6290 4 net6
rlabel metal2 s 2622 9656 2622 9656 4 net7
rlabel metal1 s 5658 10132 5658 10132 4 net8
rlabel metal1 s 3312 8398 3312 8398 4 net9
rlabel metal3 s 7199 9588 7199 9588 4 rst
flabel metal4 s 11248 496 11568 11472 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 8534 496 8854 11472 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 5820 496 6140 11472 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 3106 496 3426 11472 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 9891 496 10211 11472 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 7177 496 7497 11472 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 4463 496 4783 11472 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 1749 496 2069 11472 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 11600 5720 12000 5840 0 FreeSans 600 0 0 0 clk
port 3 nsew
flabel metal2 s 9770 11600 9826 12000 0 FreeSans 280 90 0 0 count[0]
port 4 nsew
flabel metal2 s 8482 11600 8538 12000 0 FreeSans 280 90 0 0 count[1]
port 5 nsew
flabel metal2 s 7194 11600 7250 12000 0 FreeSans 280 90 0 0 count[2]
port 6 nsew
flabel metal2 s 5906 11600 5962 12000 0 FreeSans 280 90 0 0 count[3]
port 7 nsew
flabel metal2 s 4618 11600 4674 12000 0 FreeSans 280 90 0 0 count[4]
port 8 nsew
flabel metal2 s 3330 11600 3386 12000 0 FreeSans 280 90 0 0 count[5]
port 9 nsew
flabel metal2 s 2042 11600 2098 12000 0 FreeSans 280 90 0 0 count[6]
port 10 nsew
flabel metal2 s 754 11600 810 12000 0 FreeSans 280 90 0 0 count[7]
port 11 nsew
flabel metal2 s 11058 11600 11114 12000 0 FreeSans 280 90 0 0 n_rst
port 12 nsew
<< properties >>
string FIXED_BBOX 0 0 12000 12000
string GDS_END 487306
string GDS_FILE ../gds/osc_counter.gds
string GDS_START 152836
<< end >>
