magic
tech sky130A
magscale 1 2
timestamp 1715689039
<< pwell >>
rect -201 -860 201 860
<< psubdiff >>
rect -165 790 -69 824
rect 69 790 165 824
rect -165 728 -131 790
rect 131 728 165 790
rect -165 -790 -131 -728
rect 131 -790 165 -728
rect -165 -824 -69 -790
rect 69 -824 165 -790
<< psubdiffcont >>
rect -69 790 69 824
rect -165 -728 -131 728
rect 131 -728 165 728
rect -69 -824 69 -790
<< xpolycontact >>
rect -35 262 35 694
rect -35 -694 35 -262
<< xpolyres >>
rect -35 -262 35 262
<< locali >>
rect -165 790 -69 824
rect 69 790 165 824
rect -165 728 -131 790
rect 131 728 165 790
rect -165 -790 -131 -728
rect 131 -790 165 -728
rect -165 -824 -69 -790
rect 69 -824 165 -790
<< viali >>
rect -19 279 19 676
rect -19 -676 19 -279
<< metal1 >>
rect -25 676 25 688
rect -25 279 -19 676
rect 19 279 25 676
rect -25 267 25 279
rect -25 -279 25 -267
rect -25 -676 -19 -279
rect 19 -676 25 -279
rect -25 -688 25 -676
<< properties >>
string FIXED_BBOX -148 -807 148 807
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 2.62 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 16.046k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
