magic
tech sky130A
magscale 1 2
timestamp 1715696023
<< psubdiff >>
rect -456 3854 2 3878
rect -456 3292 2 3316
<< psubdiffcont >>
rect -456 3316 2 3854
<< locali >>
rect -456 3854 2 3870
rect -456 3300 2 3316
<< viali >>
rect 4670 6266 5102 6336
rect 6398 5602 6830 5672
rect 898 5008 1330 5078
rect 2626 4344 3058 4414
rect -456 3376 2 3774
<< metal1 >>
rect 4642 6342 5128 6352
rect 4298 6336 5128 6342
rect 4298 6266 4670 6336
rect 5102 6266 5128 6336
rect 4298 6206 5128 6266
rect -768 5116 -314 5298
rect 4298 5122 4434 6206
rect 4642 6202 5128 6206
rect 6225 5672 7308 5715
rect 6225 5602 6398 5672
rect 6830 5602 7308 5672
rect 6225 5568 7308 5602
rect 7161 5123 7308 5568
rect 7806 5163 8260 5434
rect 7770 5123 8260 5163
rect -768 5078 1460 5116
rect -768 5008 898 5078
rect 1330 5008 1460 5078
rect -768 4968 1460 5008
rect 3450 4986 4454 5122
rect -768 4796 -314 4968
rect 376 3938 524 4968
rect 3450 4436 3586 4986
rect 7158 4971 8260 5123
rect 7778 4932 8260 4971
rect 2504 4414 3766 4436
rect 2504 4344 2626 4414
rect 3058 4344 3766 4414
rect 2504 4300 3766 4344
rect 3902 4300 3908 4436
rect 7778 3952 7967 4932
rect -486 3774 42 3854
rect 376 3790 1988 3938
rect -486 3376 -456 3774
rect 2 3376 42 3774
rect -486 3242 42 3376
rect -660 2760 42 3242
rect -660 2740 -206 2760
rect -562 409 -324 2740
rect -562 171 697 409
rect 935 171 941 409
rect -562 -3556 -324 171
rect -216 170 400 171
rect 1842 106 1986 3790
rect 7762 3184 7982 3952
rect 7756 2964 7762 3184
rect 7982 2964 7988 3184
rect 836 -38 842 106
rect 986 -38 1986 106
rect 7300 -3540 7484 -3534
rect -562 -3707 1883 -3556
rect 7050 -3564 7300 -3540
rect -562 -3751 -324 -3707
rect 6420 -3720 7300 -3564
rect 7050 -3724 7300 -3720
rect 7300 -3730 7484 -3724
<< via1 >>
rect 3766 4300 3902 4436
rect 697 171 935 409
rect 7762 2964 7982 3184
rect 842 -38 986 106
rect 7300 -3724 7484 -3540
<< metal2 >>
rect 3766 4436 3902 4442
rect 3766 4220 3902 4300
rect 3766 4075 3902 4084
rect 7762 3184 7982 3190
rect 7762 2481 7982 2964
rect 7758 2271 7767 2481
rect 7977 2271 7986 2481
rect 7762 2266 7982 2271
rect 697 409 935 415
rect 935 171 1065 409
rect 1303 171 1312 409
rect 697 165 935 171
rect -104 106 40 115
rect 842 106 986 112
rect 40 -38 842 106
rect -104 -47 40 -38
rect 842 -44 986 -38
rect 7294 -3724 7300 -3540
rect 7484 -3545 7638 -3540
rect 7633 -3719 7642 -3545
rect 7484 -3724 7638 -3719
<< via2 >>
rect 3766 4084 3902 4220
rect 7767 2271 7977 2481
rect 1065 171 1303 409
rect -104 -38 40 106
rect 7459 -3719 7484 -3545
rect 7484 -3719 7633 -3545
<< metal3 >>
rect 3761 4220 3907 4225
rect 3761 4084 3766 4220
rect 3902 4084 3907 4220
rect 3761 4079 3907 4084
rect 3766 4062 3902 4079
rect 3766 3920 3902 3926
rect 7762 2481 7982 2486
rect 7762 2271 7767 2481
rect 7977 2271 7982 2481
rect 1060 409 1308 414
rect 1060 171 1065 409
rect 1303 171 1373 409
rect 1611 171 1617 409
rect 1060 166 1308 171
rect 7762 159 7982 2271
rect -109 106 45 111
rect -109 -38 -104 106
rect 40 -38 45 106
rect -109 -43 45 -38
rect -104 -660 40 -43
rect 7757 -59 7763 159
rect 7981 -59 7987 159
rect 7762 -60 7982 -59
rect -104 -810 40 -804
rect 7454 -3427 7638 -3426
rect 7449 -3609 7455 -3427
rect 7637 -3609 7643 -3427
rect 7454 -3719 7459 -3609
rect 7633 -3719 7638 -3609
rect 7454 -3724 7638 -3719
<< via3 >>
rect 3766 3926 3902 4062
rect 1373 171 1611 409
rect 7763 -59 7981 159
rect -104 -804 40 -660
rect 7455 -3545 7637 -3427
rect 7455 -3609 7459 -3545
rect 7459 -3609 7633 -3545
rect 7633 -3609 7637 -3545
<< metal4 >>
rect 3765 4062 3903 4063
rect 3765 3964 3766 4062
rect 3542 3926 3766 3964
rect 3902 3964 3903 4062
rect 3902 3926 7536 3964
rect 3542 3728 7536 3926
rect 3542 2560 3778 3728
rect 7300 2448 7536 3728
rect 1716 417 1942 1932
rect 5715 417 5941 2223
rect 1372 409 1612 410
rect 1716 409 5941 417
rect 1372 171 1373 409
rect 1611 191 5941 409
rect 1611 171 1901 191
rect 1372 170 1612 171
rect 7334 159 7982 160
rect 7334 -59 7763 159
rect 7981 -59 7982 159
rect 7334 -60 7982 -59
rect -105 -660 41 -659
rect -105 -804 -104 -660
rect 40 -804 1028 -660
rect -105 -805 41 -804
rect 3564 -1158 4616 -196
rect 7334 -1028 7554 -60
rect 3820 -3282 4004 -1158
rect 3820 -3427 7638 -3282
rect 3820 -3466 7455 -3427
rect 7454 -3609 7455 -3466
rect 7637 -3609 7638 -3427
rect 7454 -3610 7638 -3609
use sky130_fd_pr__res_high_po_0p35_EMSEB3  sky130_fd_pr__res_high_po_0p35_EMSEB3_0
timestamp 1715688561
transform 0 1 5750 -1 0 5969
box -533 -1246 533 1246
use sky130_fd_pr__res_high_po_0p35_EMSEB3  sky130_fd_pr__res_high_po_0p35_EMSEB3_2
timestamp 1715688561
transform 0 1 1978 -1 0 4711
box -533 -1246 533 1246
use sky130_fd_pr__cap_mim_m3_1_MRZGNS  XC1
timestamp 1715687893
transform 1 0 2044 0 1 2192
box -1686 -1540 1686 1540
use sky130_fd_pr__cap_mim_m3_1_MRZGNS  XC2
timestamp 1715687893
transform 1 0 5784 0 1 2050
box -1686 -1540 1686 1540
use sky130_fd_pr__cap_mim_m3_1_MRZGNS  XC3
timestamp 1715687893
transform 1 0 2026 0 1 -1632
box -1686 -1540 1686 1540
use sky130_fd_pr__cap_mim_m3_1_MRZGNS  XC4
timestamp 1715687893
transform 1 0 5818 0 1 -1592
box -1686 -1540 1686 1540
use sky130_fd_pr__res_high_po_0p35_4P6F7P  XR6
timestamp 1715687893
transform 0 1 4154 -1 0 -3637
box -201 -2898 201 2898
<< labels >>
flabel metal1 -616 2860 -416 3060 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 -626 5012 -426 5212 0 FreeSans 256 0 0 0 in
port 3 nsew
flabel space 3450 4986 4704 5122 0 FreeSans 1600 0 0 0 c1_c2
flabel metal1 7902 5004 8102 5204 0 FreeSans 256 0 0 0 out
port 2 nsew
flabel metal4 3564 -1158 4616 -196 0 FreeSans 1600 0 0 0 c3_c4
<< end >>
