magic
tech sky130A
magscale 1 2
timestamp 1715770502
<< metal1 >>
rect 20418 18377 21092 18582
rect 29380 18400 30480 18860
rect 29400 18380 29880 18400
rect 20418 18272 20623 18377
rect 20412 18067 20418 18272
rect 20623 18067 20629 18272
rect 19800 16350 21150 16650
rect 20956 8129 21194 9925
rect 22150 9050 22450 9056
rect 22450 8750 25550 9050
rect 22150 8744 22450 8750
rect 20956 7891 23119 8129
rect 20956 4319 21194 7891
rect 23770 7740 23910 8750
rect 30020 8500 30480 18400
rect 29060 8040 30532 8500
rect 20956 4090 25919 4319
rect 20956 4081 23590 4090
rect 24390 4081 25919 4090
rect 22970 4080 23120 4081
rect 22970 3420 23930 3660
rect 23330 2970 23570 3420
rect 30050 2970 30290 2976
rect 23330 2730 30050 2970
rect 30050 2724 30290 2730
<< via1 >>
rect 20418 18067 20623 18272
rect 22150 8750 22450 9050
rect 30050 2730 30290 2970
<< metal2 >>
rect 20418 18272 20623 18278
rect 20418 17887 20623 18067
rect 20414 17692 20423 17887
rect 20618 17692 20627 17887
rect 20418 17687 20623 17692
rect 19656 8750 22150 9050
rect 22450 8750 22456 9050
rect 25850 5530 26090 5550
rect 25850 5420 25870 5530
rect 25990 5420 26090 5530
rect 25850 5260 26090 5420
rect 27920 5430 28180 5450
rect 27920 5290 28040 5430
rect 28160 5290 28180 5430
rect 27920 5250 28180 5290
rect 30050 4420 30290 4429
rect 30050 2970 30290 4180
rect 30044 2730 30050 2970
rect 30290 2730 30296 2970
<< via2 >>
rect 20423 17692 20618 17887
rect 25870 5420 25990 5530
rect 28040 5290 28160 5430
rect 30050 4180 30290 4420
<< metal3 >>
rect 20418 17887 20623 17892
rect 20418 17692 20423 17887
rect 20618 17692 20623 17887
rect 20418 5500 20623 17692
rect 24660 5530 26030 5570
rect 24660 5500 25870 5530
rect 20418 5420 25870 5500
rect 25990 5420 26030 5530
rect 20418 5390 26030 5420
rect 28030 5460 30000 5480
rect 28030 5430 30290 5460
rect 20418 5300 24790 5390
rect 20418 5298 20623 5300
rect 28030 5290 28040 5430
rect 28160 5320 30290 5430
rect 28160 5290 28190 5320
rect 28030 5280 28190 5290
rect 29830 5220 30290 5320
rect 30050 4425 30290 5220
rect 30045 4420 30295 4425
rect 30045 4180 30050 4420
rect 30290 4180 30295 4420
rect 30045 4175 30295 4180
use p3_opamp  p3_opamp_0
timestamp 1715689418
transform 1 0 21230 0 1 920
box 3650 3170 8500 8260
use sky130_fd_pr__res_high_po_0p35_5FS976  sky130_fd_pr__res_high_po_0p35_5FS976_0
timestamp 1715691009
transform -1 0 23851 0 -1 5768
box -201 -2598 201 2598
use sky130_fd_pr__res_high_po_0p35_5FS976  sky130_fd_pr__res_high_po_0p35_5FS976_1
timestamp 1715691009
transform 1 0 23041 0 1 5728
box -201 -2598 201 2598
use twin_tee  twin_tee_0
timestamp 1715696023
transform 1 0 21518 0 1 13438
box -768 -3838 8260 6502
<< labels >>
flabel metal1 19800 16350 21150 16650 0 FreeSans 1600 0 0 0 vss
port 1 nsew
flabel metal2 19656 8750 22150 9050 0 FreeSans 1600 0 0 0 vdd
port 2 nsew
flabel metal1 30020 8040 30480 18860 0 FreeSans 1600 0 0 0 out
port 4 nsew
<< properties >>
<< end >>
