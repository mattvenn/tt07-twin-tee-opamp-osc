magic
tech sky130A
magscale 1 2
timestamp 1715687893
<< metal3 >>
rect -1686 1512 1686 1540
rect -1686 -1512 1602 1512
rect 1666 -1512 1686 1512
rect -1686 -1540 1686 -1512
<< via3 >>
rect 1602 -1512 1666 1512
<< mimcap >>
rect -1646 1460 1354 1500
rect -1646 -1460 -1606 1460
rect 1314 -1460 1354 1460
rect -1646 -1500 1354 -1460
<< mimcapcontact >>
rect -1606 -1460 1314 1460
<< metal4 >>
rect 1586 1512 1682 1528
rect -1607 1460 1315 1461
rect -1607 -1460 -1606 1460
rect 1314 -1460 1315 1460
rect -1607 -1461 1315 -1460
rect 1586 -1512 1602 1512
rect 1666 -1512 1682 1512
rect 1586 -1528 1682 -1512
<< properties >>
string FIXED_BBOX -1686 -1540 1394 1540
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 15.0 l 15.0 val 461.4 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
