VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_twin_tee_opamp_osc
  CLASS BLOCK ;
  FOREIGN tt_um_twin_tee_opamp_osc ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.060000 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 130.800 94.380 143.260 99.710 ;
        RECT 111.940 88.090 124.400 93.420 ;
        RECT 114.560 48.010 143.540 50.020 ;
        RECT 114.890 15.660 116.900 41.640 ;
        RECT 118.940 15.860 120.950 41.840 ;
        RECT 126.840 34.010 128.850 42.890 ;
        RECT 126.290 22.360 129.390 33.190 ;
      LAYER nwell ;
        RECT 130.890 28.410 134.080 43.820 ;
        RECT 137.240 28.410 140.430 43.820 ;
      LAYER pwell ;
        RECT 131.040 25.560 140.240 28.020 ;
      LAYER nwell ;
        RECT 141.840 26.610 145.030 44.080 ;
      LAYER pwell ;
        RECT 137.840 25.510 138.390 25.560 ;
        RECT 130.340 22.410 141.170 25.510 ;
        RECT 145.840 22.410 148.940 40.110 ;
      LAYER li1 ;
        RECT 130.980 99.360 143.080 99.530 ;
        RECT 130.980 94.730 131.150 99.360 ;
        RECT 131.630 98.530 133.790 98.880 ;
        RECT 140.270 95.210 142.430 95.560 ;
        RECT 142.910 94.730 143.080 99.360 ;
        RECT 130.980 94.560 143.080 94.730 ;
        RECT 112.120 93.070 124.220 93.240 ;
        RECT 112.120 88.440 112.290 93.070 ;
        RECT 112.770 92.240 114.930 92.590 ;
        RECT 121.410 88.920 123.570 89.270 ;
        RECT 124.050 88.440 124.220 93.070 ;
        RECT 112.120 88.270 124.220 88.440 ;
        RECT 106.000 83.700 108.290 86.550 ;
        RECT 114.740 49.670 143.360 49.840 ;
        RECT 114.740 48.360 114.910 49.670 ;
        RECT 115.390 48.840 117.550 49.190 ;
        RECT 140.550 48.840 142.710 49.190 ;
        RECT 143.190 48.360 143.360 49.670 ;
        RECT 114.740 48.190 143.360 48.360 ;
        RECT 142.020 43.730 144.850 43.900 ;
        RECT 131.070 43.470 133.900 43.640 ;
        RECT 131.070 43.110 131.240 43.470 ;
        RECT 127.020 42.540 128.670 42.710 ;
        RECT 127.020 42.410 127.190 42.540 ;
        RECT 119.120 41.490 120.770 41.660 ;
        RECT 115.070 41.290 116.720 41.460 ;
        RECT 115.070 16.010 115.240 41.290 ;
        RECT 115.720 38.650 116.070 40.810 ;
        RECT 115.720 16.490 116.070 18.650 ;
        RECT 116.550 16.010 116.720 41.290 ;
        RECT 119.120 16.210 119.290 41.490 ;
        RECT 119.770 38.850 120.120 41.010 ;
        RECT 119.770 16.690 120.120 18.850 ;
        RECT 120.600 16.210 120.770 41.490 ;
        RECT 125.190 34.360 127.190 42.410 ;
        RECT 127.670 39.900 128.020 42.060 ;
        RECT 127.670 34.840 128.020 37.000 ;
        RECT 128.500 34.360 128.670 42.540 ;
        RECT 125.190 34.190 128.670 34.360 ;
        RECT 125.190 33.010 128.340 34.190 ;
        RECT 125.190 32.840 129.210 33.010 ;
        RECT 125.190 22.710 126.640 32.840 ;
        RECT 127.320 32.270 128.360 32.440 ;
        RECT 126.980 30.210 127.150 32.210 ;
        RECT 128.530 30.210 128.700 32.210 ;
        RECT 127.320 29.980 128.360 30.150 ;
        RECT 126.980 27.920 127.150 29.920 ;
        RECT 128.530 27.920 128.700 29.920 ;
        RECT 127.320 27.690 128.360 27.860 ;
        RECT 126.980 25.630 127.150 27.630 ;
        RECT 128.530 25.630 128.700 27.630 ;
        RECT 127.320 25.400 128.360 25.570 ;
        RECT 126.980 23.340 127.150 25.340 ;
        RECT 128.530 23.340 128.700 25.340 ;
        RECT 129.040 25.010 129.210 32.840 ;
        RECT 130.940 31.210 131.240 43.110 ;
        RECT 131.965 42.900 133.005 43.070 ;
        RECT 131.580 40.840 131.750 42.840 ;
        RECT 133.220 40.840 133.390 42.840 ;
        RECT 131.965 40.610 133.005 40.780 ;
        RECT 131.580 38.550 131.750 40.550 ;
        RECT 133.220 38.550 133.390 40.550 ;
        RECT 131.965 38.320 133.005 38.490 ;
        RECT 131.580 36.260 131.750 38.260 ;
        RECT 133.220 36.260 133.390 38.260 ;
        RECT 131.965 36.030 133.005 36.200 ;
        RECT 131.580 33.970 131.750 35.970 ;
        RECT 133.220 33.970 133.390 35.970 ;
        RECT 131.965 33.740 133.005 33.910 ;
        RECT 131.580 31.680 131.750 33.680 ;
        RECT 133.220 31.680 133.390 33.680 ;
        RECT 131.965 31.450 133.005 31.620 ;
        RECT 131.070 28.760 131.240 31.210 ;
        RECT 131.580 29.390 131.750 31.390 ;
        RECT 133.220 29.390 133.390 31.390 ;
        RECT 131.965 29.160 133.005 29.330 ;
        RECT 133.730 28.760 133.900 43.470 ;
        RECT 131.070 28.590 133.900 28.760 ;
        RECT 137.420 43.470 140.250 43.640 ;
        RECT 137.420 28.760 137.590 43.470 ;
        RECT 140.080 43.110 140.250 43.470 ;
        RECT 142.020 43.360 142.190 43.730 ;
        RECT 138.315 42.900 139.355 43.070 ;
        RECT 137.930 40.840 138.100 42.840 ;
        RECT 139.570 40.840 139.740 42.840 ;
        RECT 138.315 40.610 139.355 40.780 ;
        RECT 137.930 38.550 138.100 40.550 ;
        RECT 139.570 38.550 139.740 40.550 ;
        RECT 138.315 38.320 139.355 38.490 ;
        RECT 137.930 36.260 138.100 38.260 ;
        RECT 139.570 36.260 139.740 38.260 ;
        RECT 138.315 36.030 139.355 36.200 ;
        RECT 137.930 33.970 138.100 35.970 ;
        RECT 139.570 33.970 139.740 35.970 ;
        RECT 138.315 33.740 139.355 33.910 ;
        RECT 137.930 31.680 138.100 33.680 ;
        RECT 139.570 31.680 139.740 33.680 ;
        RECT 138.315 31.450 139.355 31.620 ;
        RECT 137.930 29.390 138.100 31.390 ;
        RECT 139.570 29.390 139.740 31.390 ;
        RECT 140.080 31.210 140.390 43.110 ;
        RECT 138.315 29.160 139.355 29.330 ;
        RECT 140.080 28.760 140.250 31.210 ;
        RECT 137.420 28.590 140.250 28.760 ;
        RECT 131.220 27.670 135.460 27.840 ;
        RECT 131.220 25.910 131.390 27.670 ;
        RECT 132.070 27.100 134.610 27.270 ;
        RECT 131.730 26.540 131.900 27.040 ;
        RECT 134.780 26.540 134.950 27.040 ;
        RECT 132.070 26.310 134.610 26.480 ;
        RECT 135.290 25.910 135.460 27.670 ;
        RECT 131.220 25.740 135.460 25.910 ;
        RECT 135.820 27.670 140.060 27.840 ;
        RECT 141.990 27.810 142.190 43.360 ;
        RECT 142.915 43.160 143.955 43.330 ;
        RECT 142.530 42.600 142.700 43.100 ;
        RECT 144.170 42.600 144.340 43.100 ;
        RECT 142.915 42.370 143.955 42.540 ;
        RECT 142.530 41.810 142.700 42.310 ;
        RECT 144.170 41.810 144.340 42.310 ;
        RECT 142.915 41.580 143.955 41.750 ;
        RECT 142.530 41.020 142.700 41.520 ;
        RECT 144.170 41.020 144.340 41.520 ;
        RECT 142.915 40.790 143.955 40.960 ;
        RECT 142.530 40.230 142.700 40.730 ;
        RECT 144.170 40.230 144.340 40.730 ;
        RECT 142.915 40.000 143.955 40.170 ;
        RECT 142.530 39.440 142.700 39.940 ;
        RECT 144.170 39.440 144.340 39.940 ;
        RECT 142.915 39.210 143.955 39.380 ;
        RECT 142.530 38.650 142.700 39.150 ;
        RECT 144.170 38.650 144.340 39.150 ;
        RECT 142.915 38.420 143.955 38.590 ;
        RECT 142.530 37.860 142.700 38.360 ;
        RECT 144.170 37.860 144.340 38.360 ;
        RECT 142.915 37.630 143.955 37.800 ;
        RECT 142.530 37.070 142.700 37.570 ;
        RECT 144.170 37.070 144.340 37.570 ;
        RECT 142.915 36.840 143.955 37.010 ;
        RECT 142.530 36.280 142.700 36.780 ;
        RECT 144.170 36.280 144.340 36.780 ;
        RECT 142.915 36.050 143.955 36.220 ;
        RECT 142.530 35.490 142.700 35.990 ;
        RECT 144.170 35.490 144.340 35.990 ;
        RECT 142.915 35.260 143.955 35.430 ;
        RECT 142.530 34.700 142.700 35.200 ;
        RECT 144.170 34.700 144.340 35.200 ;
        RECT 142.915 34.470 143.955 34.640 ;
        RECT 142.530 33.910 142.700 34.410 ;
        RECT 144.170 33.910 144.340 34.410 ;
        RECT 142.915 33.680 143.955 33.850 ;
        RECT 142.530 33.120 142.700 33.620 ;
        RECT 144.170 33.120 144.340 33.620 ;
        RECT 142.915 32.890 143.955 33.060 ;
        RECT 142.530 32.330 142.700 32.830 ;
        RECT 144.170 32.330 144.340 32.830 ;
        RECT 142.915 32.100 143.955 32.270 ;
        RECT 142.530 31.540 142.700 32.040 ;
        RECT 144.170 31.540 144.340 32.040 ;
        RECT 142.915 31.310 143.955 31.480 ;
        RECT 142.530 30.750 142.700 31.250 ;
        RECT 144.170 30.750 144.340 31.250 ;
        RECT 142.915 30.520 143.955 30.690 ;
        RECT 142.530 29.960 142.700 30.460 ;
        RECT 144.170 29.960 144.340 30.460 ;
        RECT 142.915 29.730 143.955 29.900 ;
        RECT 142.530 29.170 142.700 29.670 ;
        RECT 144.170 29.170 144.340 29.670 ;
        RECT 142.915 28.940 143.955 29.110 ;
        RECT 142.530 28.380 142.700 28.880 ;
        RECT 144.170 28.380 144.340 28.880 ;
        RECT 142.915 28.150 143.955 28.320 ;
        RECT 135.820 25.910 135.990 27.670 ;
        RECT 136.670 27.100 139.210 27.270 ;
        RECT 136.330 26.540 136.500 27.040 ;
        RECT 139.380 26.540 139.550 27.040 ;
        RECT 136.670 26.310 139.210 26.480 ;
        RECT 139.890 25.910 140.060 27.670 ;
        RECT 142.020 26.960 142.190 27.810 ;
        RECT 142.530 27.590 142.700 28.090 ;
        RECT 144.170 27.590 144.340 28.090 ;
        RECT 142.915 27.360 143.955 27.530 ;
        RECT 144.680 26.960 144.850 43.730 ;
        RECT 142.020 26.790 144.850 26.960 ;
        RECT 146.020 39.760 148.760 39.930 ;
        RECT 135.820 25.740 140.190 25.910 ;
        RECT 131.240 25.710 132.040 25.740 ;
        RECT 139.390 25.710 140.190 25.740 ;
        RECT 130.520 25.260 140.990 25.330 ;
        RECT 146.020 25.260 146.190 39.760 ;
        RECT 146.870 39.190 147.910 39.360 ;
        RECT 146.530 37.130 146.700 39.130 ;
        RECT 148.080 37.130 148.250 39.130 ;
        RECT 146.870 36.900 147.910 37.070 ;
        RECT 148.590 37.060 148.760 39.760 ;
        RECT 146.530 34.840 146.700 36.840 ;
        RECT 148.080 34.840 148.250 36.840 ;
        RECT 146.870 34.610 147.910 34.780 ;
        RECT 146.530 32.550 146.700 34.550 ;
        RECT 148.080 32.550 148.250 34.550 ;
        RECT 146.870 32.320 147.910 32.490 ;
        RECT 146.530 30.260 146.700 32.260 ;
        RECT 148.080 30.260 148.250 32.260 ;
        RECT 146.870 30.030 147.910 30.200 ;
        RECT 146.530 27.970 146.700 29.970 ;
        RECT 148.080 27.970 148.250 29.970 ;
        RECT 146.870 27.740 147.910 27.910 ;
        RECT 146.530 25.680 146.700 27.680 ;
        RECT 148.080 25.680 148.250 27.680 ;
        RECT 146.870 25.450 147.910 25.620 ;
        RECT 130.520 25.160 146.190 25.260 ;
        RECT 130.520 25.010 130.690 25.160 ;
        RECT 127.320 23.110 128.360 23.280 ;
        RECT 129.040 22.760 130.690 25.010 ;
        RECT 131.320 24.650 133.320 24.820 ;
        RECT 133.610 24.650 135.610 24.820 ;
        RECT 135.900 24.650 137.900 24.820 ;
        RECT 138.190 24.650 140.190 24.820 ;
        RECT 140.820 24.660 146.190 25.160 ;
        RECT 131.090 23.440 131.260 24.480 ;
        RECT 133.380 23.440 133.550 24.480 ;
        RECT 135.670 23.440 135.840 24.480 ;
        RECT 137.960 23.440 138.130 24.480 ;
        RECT 140.250 23.440 140.420 24.480 ;
        RECT 131.320 23.100 133.320 23.270 ;
        RECT 133.610 23.100 135.610 23.270 ;
        RECT 135.900 23.100 137.900 23.270 ;
        RECT 138.190 23.100 140.190 23.270 ;
        RECT 140.790 23.060 146.190 24.660 ;
        RECT 146.530 23.390 146.700 25.390 ;
        RECT 148.080 23.390 148.250 25.390 ;
        RECT 146.870 23.160 147.910 23.330 ;
        RECT 140.820 22.760 146.190 23.060 ;
        RECT 148.590 22.760 149.340 37.060 ;
        RECT 126.890 22.710 128.790 22.760 ;
        RECT 129.040 22.710 149.340 22.760 ;
        RECT 125.190 20.510 149.340 22.710 ;
        RECT 119.120 16.040 120.770 16.210 ;
        RECT 115.070 15.840 116.720 16.010 ;
      LAYER mcon ;
        RECT 106.000 84.080 108.290 86.070 ;
        RECT 115.480 48.920 117.465 49.110 ;
        RECT 140.635 48.920 142.620 49.110 ;
        RECT 115.800 38.735 115.990 40.720 ;
        RECT 115.800 16.580 115.990 18.565 ;
        RECT 119.850 38.935 120.040 40.920 ;
        RECT 119.850 16.780 120.040 18.765 ;
        RECT 125.690 38.110 126.540 41.810 ;
        RECT 126.940 34.810 127.190 41.960 ;
        RECT 127.750 39.985 127.940 41.970 ;
        RECT 127.750 34.930 127.940 36.915 ;
        RECT 126.390 23.560 126.640 32.910 ;
        RECT 127.400 32.270 128.280 32.440 ;
        RECT 126.980 30.290 127.150 32.130 ;
        RECT 128.530 30.290 128.700 32.130 ;
        RECT 127.400 29.980 128.280 30.150 ;
        RECT 126.980 28.000 127.150 29.840 ;
        RECT 128.530 28.000 128.700 29.840 ;
        RECT 127.400 27.690 128.280 27.860 ;
        RECT 126.980 25.710 127.150 27.550 ;
        RECT 128.530 25.710 128.700 27.550 ;
        RECT 127.400 25.400 128.280 25.570 ;
        RECT 126.980 23.420 127.150 25.260 ;
        RECT 128.530 23.420 128.700 25.260 ;
        RECT 130.940 31.210 131.240 43.110 ;
        RECT 132.045 42.900 132.925 43.070 ;
        RECT 131.580 40.920 131.750 42.760 ;
        RECT 133.220 40.920 133.390 42.760 ;
        RECT 132.045 40.610 132.925 40.780 ;
        RECT 131.580 38.630 131.750 40.470 ;
        RECT 133.220 38.630 133.390 40.470 ;
        RECT 132.045 38.320 132.925 38.490 ;
        RECT 131.580 36.340 131.750 38.180 ;
        RECT 133.220 36.340 133.390 38.180 ;
        RECT 132.045 36.030 132.925 36.200 ;
        RECT 131.580 34.050 131.750 35.890 ;
        RECT 133.220 34.050 133.390 35.890 ;
        RECT 132.045 33.740 132.925 33.910 ;
        RECT 131.580 31.760 131.750 33.600 ;
        RECT 133.220 31.760 133.390 33.600 ;
        RECT 132.045 31.450 132.925 31.620 ;
        RECT 131.580 29.470 131.750 31.310 ;
        RECT 133.220 29.470 133.390 31.310 ;
        RECT 132.045 29.160 132.925 29.330 ;
        RECT 138.395 42.900 139.275 43.070 ;
        RECT 137.930 40.920 138.100 42.760 ;
        RECT 139.570 40.920 139.740 42.760 ;
        RECT 138.395 40.610 139.275 40.780 ;
        RECT 137.930 38.630 138.100 40.470 ;
        RECT 139.570 38.630 139.740 40.470 ;
        RECT 138.395 38.320 139.275 38.490 ;
        RECT 137.930 36.340 138.100 38.180 ;
        RECT 139.570 36.340 139.740 38.180 ;
        RECT 138.395 36.030 139.275 36.200 ;
        RECT 137.930 34.050 138.100 35.890 ;
        RECT 139.570 34.050 139.740 35.890 ;
        RECT 138.395 33.740 139.275 33.910 ;
        RECT 137.930 31.760 138.100 33.600 ;
        RECT 139.570 31.760 139.740 33.600 ;
        RECT 138.395 31.450 139.275 31.620 ;
        RECT 137.930 29.470 138.100 31.310 ;
        RECT 139.570 29.470 139.740 31.310 ;
        RECT 140.090 31.210 140.390 43.110 ;
        RECT 138.395 29.160 139.275 29.330 ;
        RECT 132.150 27.100 134.530 27.270 ;
        RECT 131.730 26.620 131.900 26.960 ;
        RECT 134.780 26.620 134.950 26.960 ;
        RECT 132.150 26.310 134.530 26.480 ;
        RECT 141.990 27.810 142.190 43.360 ;
        RECT 142.995 43.160 143.875 43.330 ;
        RECT 142.530 42.680 142.700 43.020 ;
        RECT 144.170 42.680 144.340 43.020 ;
        RECT 142.995 42.370 143.875 42.540 ;
        RECT 142.530 41.890 142.700 42.230 ;
        RECT 144.170 41.890 144.340 42.230 ;
        RECT 142.995 41.580 143.875 41.750 ;
        RECT 142.530 41.100 142.700 41.440 ;
        RECT 144.170 41.100 144.340 41.440 ;
        RECT 142.995 40.790 143.875 40.960 ;
        RECT 142.530 40.310 142.700 40.650 ;
        RECT 144.170 40.310 144.340 40.650 ;
        RECT 142.995 40.000 143.875 40.170 ;
        RECT 142.530 39.520 142.700 39.860 ;
        RECT 144.170 39.520 144.340 39.860 ;
        RECT 142.995 39.210 143.875 39.380 ;
        RECT 142.530 38.730 142.700 39.070 ;
        RECT 144.170 38.730 144.340 39.070 ;
        RECT 142.995 38.420 143.875 38.590 ;
        RECT 142.530 37.940 142.700 38.280 ;
        RECT 144.170 37.940 144.340 38.280 ;
        RECT 142.995 37.630 143.875 37.800 ;
        RECT 142.530 37.150 142.700 37.490 ;
        RECT 144.170 37.150 144.340 37.490 ;
        RECT 142.995 36.840 143.875 37.010 ;
        RECT 142.530 36.360 142.700 36.700 ;
        RECT 144.170 36.360 144.340 36.700 ;
        RECT 142.995 36.050 143.875 36.220 ;
        RECT 142.530 35.570 142.700 35.910 ;
        RECT 144.170 35.570 144.340 35.910 ;
        RECT 142.995 35.260 143.875 35.430 ;
        RECT 142.530 34.780 142.700 35.120 ;
        RECT 144.170 34.780 144.340 35.120 ;
        RECT 142.995 34.470 143.875 34.640 ;
        RECT 142.530 33.990 142.700 34.330 ;
        RECT 144.170 33.990 144.340 34.330 ;
        RECT 142.995 33.680 143.875 33.850 ;
        RECT 142.530 33.200 142.700 33.540 ;
        RECT 144.170 33.200 144.340 33.540 ;
        RECT 142.995 32.890 143.875 33.060 ;
        RECT 142.530 32.410 142.700 32.750 ;
        RECT 144.170 32.410 144.340 32.750 ;
        RECT 142.995 32.100 143.875 32.270 ;
        RECT 142.530 31.620 142.700 31.960 ;
        RECT 144.170 31.620 144.340 31.960 ;
        RECT 142.995 31.310 143.875 31.480 ;
        RECT 142.530 30.830 142.700 31.170 ;
        RECT 144.170 30.830 144.340 31.170 ;
        RECT 142.995 30.520 143.875 30.690 ;
        RECT 142.530 30.040 142.700 30.380 ;
        RECT 144.170 30.040 144.340 30.380 ;
        RECT 142.995 29.730 143.875 29.900 ;
        RECT 142.530 29.250 142.700 29.590 ;
        RECT 144.170 29.250 144.340 29.590 ;
        RECT 142.995 28.940 143.875 29.110 ;
        RECT 142.530 28.460 142.700 28.800 ;
        RECT 144.170 28.460 144.340 28.800 ;
        RECT 142.995 28.150 143.875 28.320 ;
        RECT 136.750 27.100 139.130 27.270 ;
        RECT 136.330 26.620 136.500 26.960 ;
        RECT 139.380 26.620 139.550 26.960 ;
        RECT 136.750 26.310 139.130 26.480 ;
        RECT 142.530 27.670 142.700 28.010 ;
        RECT 144.170 27.670 144.340 28.010 ;
        RECT 142.995 27.360 143.875 27.530 ;
        RECT 146.950 39.190 147.830 39.360 ;
        RECT 146.530 37.210 146.700 39.050 ;
        RECT 148.080 37.210 148.250 39.050 ;
        RECT 146.950 36.900 147.830 37.070 ;
        RECT 146.530 34.920 146.700 36.760 ;
        RECT 148.080 34.920 148.250 36.760 ;
        RECT 146.950 34.610 147.830 34.780 ;
        RECT 146.530 32.630 146.700 34.470 ;
        RECT 148.080 32.630 148.250 34.470 ;
        RECT 146.950 32.320 147.830 32.490 ;
        RECT 146.530 30.340 146.700 32.180 ;
        RECT 148.080 30.340 148.250 32.180 ;
        RECT 146.950 30.030 147.830 30.200 ;
        RECT 146.530 28.050 146.700 29.890 ;
        RECT 148.080 28.050 148.250 29.890 ;
        RECT 146.950 27.740 147.830 27.910 ;
        RECT 146.530 25.760 146.700 27.600 ;
        RECT 148.080 25.760 148.250 27.600 ;
        RECT 146.950 25.450 147.830 25.620 ;
        RECT 127.400 23.110 128.280 23.280 ;
        RECT 131.400 24.650 133.240 24.820 ;
        RECT 133.690 24.650 135.530 24.820 ;
        RECT 135.980 24.650 137.820 24.820 ;
        RECT 138.270 24.650 140.110 24.820 ;
        RECT 131.090 23.520 131.260 24.400 ;
        RECT 133.380 23.520 133.550 24.400 ;
        RECT 135.670 23.520 135.840 24.400 ;
        RECT 137.960 23.520 138.130 24.400 ;
        RECT 140.250 23.520 140.420 24.400 ;
        RECT 131.400 23.100 133.240 23.270 ;
        RECT 133.690 23.100 135.530 23.270 ;
        RECT 135.980 23.100 137.820 23.270 ;
        RECT 138.270 23.100 140.110 23.270 ;
        RECT 145.940 23.060 146.190 24.210 ;
        RECT 146.530 23.470 146.700 25.310 ;
        RECT 148.080 23.470 148.250 25.310 ;
        RECT 146.950 23.160 147.830 23.330 ;
        RECT 148.590 23.060 148.840 24.210 ;
        RECT 126.890 22.460 128.790 22.760 ;
        RECT 130.990 22.510 140.540 22.760 ;
        RECT 146.290 22.560 148.490 22.760 ;
        RECT 128.490 20.810 147.440 21.360 ;
      LAYER met1 ;
        RECT 131.490 98.910 133.920 98.960 ;
        RECT 129.770 98.230 133.920 98.910 ;
        RECT 104.440 92.920 106.710 93.690 ;
        RECT 102.780 92.780 106.710 92.920 ;
        RECT 129.770 92.810 130.450 98.230 ;
        RECT 131.490 98.210 133.920 98.230 ;
        RECT 139.405 95.040 144.820 95.775 ;
        RECT 144.085 92.815 144.820 95.040 ;
        RECT 147.310 94.310 149.580 94.370 ;
        RECT 147.310 93.015 153.090 94.310 ;
        RECT 147.130 92.815 153.090 93.015 ;
        RECT 102.780 92.040 115.580 92.780 ;
        RECT 125.530 92.130 130.550 92.810 ;
        RECT 102.780 91.895 106.710 92.040 ;
        RECT 102.780 91.370 103.805 91.895 ;
        RECT 102.750 90.345 103.835 91.370 ;
        RECT 104.440 91.180 106.710 91.895 ;
        RECT 110.160 86.890 110.900 92.040 ;
        RECT 125.530 89.380 126.210 92.130 ;
        RECT 144.070 92.055 153.090 92.815 ;
        RECT 147.170 92.010 153.090 92.055 ;
        RECT 147.170 91.910 150.090 92.010 ;
        RECT 147.170 91.860 149.580 91.910 ;
        RECT 120.800 88.700 127.820 89.380 ;
        RECT 147.170 86.960 148.115 91.860 ;
        RECT 105.850 83.410 108.490 86.470 ;
        RECT 110.160 86.150 118.220 86.890 ;
        RECT 93.750 83.250 95.250 83.280 ;
        RECT 104.980 83.260 108.490 83.410 ;
        RECT 99.690 83.250 108.490 83.260 ;
        RECT 93.750 81.760 108.490 83.250 ;
        RECT 93.750 81.750 99.710 81.760 ;
        RECT 93.750 81.720 95.250 81.750 ;
        RECT 104.980 81.000 108.490 81.760 ;
        RECT 104.980 80.900 107.250 81.000 ;
        RECT 105.470 69.245 106.660 80.900 ;
        RECT 105.470 68.055 112.985 69.245 ;
        RECT 105.470 49.420 106.660 68.055 ;
        RECT 107.200 68.050 110.280 68.055 ;
        RECT 117.490 67.730 118.210 86.150 ;
        RECT 147.090 83.120 148.190 86.960 ;
        RECT 147.060 82.020 148.220 83.120 ;
        RECT 112.460 67.010 118.210 67.730 ;
        RECT 144.780 49.500 145.700 49.530 ;
        RECT 105.470 48.665 117.695 49.420 ;
        RECT 143.530 49.380 145.700 49.500 ;
        RECT 105.470 40.655 106.660 48.665 ;
        RECT 140.380 48.600 145.700 49.380 ;
        RECT 143.530 48.580 145.700 48.600 ;
        RECT 144.780 48.550 145.700 48.580 ;
        RECT 111.440 45.260 112.940 45.290 ;
        RECT 125.090 45.260 149.340 45.910 ;
        RECT 111.440 43.760 149.340 45.260 ;
        RECT 111.440 43.730 112.940 43.760 ;
        RECT 115.770 40.655 116.020 40.780 ;
        RECT 105.470 39.465 116.285 40.655 ;
        RECT 105.470 21.605 106.660 39.465 ;
        RECT 115.770 38.675 116.020 39.465 ;
        RECT 119.540 38.710 120.240 43.760 ;
        RECT 125.090 43.560 149.340 43.760 ;
        RECT 125.090 34.660 127.290 42.410 ;
        RECT 127.440 39.660 128.390 43.560 ;
        RECT 127.720 36.960 127.970 36.975 ;
        RECT 125.090 22.810 126.740 34.660 ;
        RECT 127.590 34.460 129.440 36.960 ;
        RECT 127.340 32.210 128.340 32.560 ;
        RECT 126.950 31.760 127.180 32.190 ;
        RECT 128.490 31.760 129.440 34.460 ;
        RECT 126.940 30.610 129.440 31.760 ;
        RECT 129.590 31.060 131.340 43.560 ;
        RECT 131.940 42.860 137.290 43.210 ;
        RECT 138.290 42.860 139.390 43.160 ;
        RECT 131.550 42.460 131.780 42.820 ;
        RECT 133.140 42.810 137.290 42.860 ;
        RECT 133.140 42.460 137.640 42.810 ;
        RECT 137.900 42.460 138.130 42.820 ;
        RECT 139.540 42.460 139.770 42.820 ;
        RECT 131.540 41.660 139.770 42.460 ;
        RECT 131.540 41.260 135.140 41.660 ;
        RECT 131.550 40.860 131.780 41.260 ;
        RECT 133.140 41.210 135.140 41.260 ;
        RECT 133.190 40.860 135.140 41.210 ;
        RECT 131.990 40.810 132.990 40.860 ;
        RECT 131.985 40.580 132.990 40.810 ;
        RECT 131.990 40.560 132.990 40.580 ;
        RECT 133.240 40.530 135.140 40.860 ;
        RECT 131.550 40.110 131.780 40.530 ;
        RECT 133.190 40.110 135.140 40.530 ;
        RECT 131.540 38.860 135.140 40.110 ;
        RECT 131.550 38.570 131.780 38.860 ;
        RECT 133.140 38.560 135.140 38.860 ;
        RECT 131.940 38.260 135.140 38.560 ;
        RECT 131.550 37.960 131.780 38.240 ;
        RECT 133.140 37.960 135.140 38.260 ;
        RECT 131.540 36.760 135.140 37.960 ;
        RECT 131.550 36.280 131.780 36.760 ;
        RECT 131.990 36.230 132.990 36.260 ;
        RECT 131.985 36.000 132.990 36.230 ;
        RECT 131.990 35.960 132.990 36.000 ;
        RECT 131.550 35.660 131.780 35.950 ;
        RECT 133.140 35.660 135.140 36.760 ;
        RECT 131.540 34.460 135.140 35.660 ;
        RECT 131.550 33.990 131.780 34.460 ;
        RECT 133.140 33.960 135.140 34.460 ;
        RECT 131.940 33.710 135.140 33.960 ;
        RECT 131.550 33.260 131.780 33.660 ;
        RECT 133.140 33.260 135.140 33.710 ;
        RECT 131.540 32.060 135.140 33.260 ;
        RECT 131.550 31.700 131.780 32.060 ;
        RECT 131.990 31.650 132.990 31.710 ;
        RECT 131.985 31.420 132.990 31.650 ;
        RECT 131.990 31.410 132.990 31.420 ;
        RECT 131.550 31.010 131.780 31.370 ;
        RECT 133.140 31.010 135.140 32.060 ;
        RECT 126.950 30.230 127.180 30.610 ;
        RECT 128.490 30.210 129.440 30.610 ;
        RECT 127.340 29.910 129.440 30.210 ;
        RECT 126.950 29.510 127.180 29.900 ;
        RECT 128.490 29.510 129.440 29.910 ;
        RECT 131.540 29.810 135.140 31.010 ;
        RECT 126.940 28.360 129.440 29.510 ;
        RECT 131.550 29.410 131.780 29.810 ;
        RECT 133.140 29.360 135.140 29.810 ;
        RECT 131.940 29.160 135.140 29.360 ;
        RECT 136.140 41.260 139.770 41.660 ;
        RECT 136.140 40.060 137.640 41.260 ;
        RECT 137.900 40.860 138.130 41.260 ;
        RECT 139.540 40.860 139.770 41.260 ;
        RECT 138.340 40.810 139.390 40.860 ;
        RECT 138.335 40.580 139.390 40.810 ;
        RECT 138.340 40.560 139.390 40.580 ;
        RECT 137.900 40.060 138.130 40.530 ;
        RECT 139.540 40.060 139.770 40.530 ;
        RECT 136.140 38.860 139.770 40.060 ;
        RECT 136.140 37.960 137.640 38.860 ;
        RECT 137.900 38.570 138.130 38.860 ;
        RECT 139.540 38.570 139.770 38.860 ;
        RECT 138.290 38.260 139.390 38.560 ;
        RECT 137.900 37.960 138.130 38.240 ;
        RECT 139.540 37.960 139.770 38.240 ;
        RECT 136.140 36.760 139.770 37.960 ;
        RECT 136.140 35.660 137.640 36.760 ;
        RECT 137.900 36.280 138.130 36.760 ;
        RECT 139.540 36.280 139.770 36.760 ;
        RECT 138.340 36.230 139.390 36.260 ;
        RECT 138.335 36.000 139.390 36.230 ;
        RECT 138.340 35.960 139.390 36.000 ;
        RECT 137.900 35.660 138.130 35.950 ;
        RECT 139.540 35.660 139.770 35.950 ;
        RECT 136.140 34.460 139.770 35.660 ;
        RECT 136.140 33.260 137.640 34.460 ;
        RECT 137.900 33.990 138.130 34.460 ;
        RECT 139.540 33.990 139.770 34.460 ;
        RECT 138.290 33.660 139.390 33.960 ;
        RECT 137.900 33.260 138.130 33.660 ;
        RECT 139.540 33.260 139.770 33.660 ;
        RECT 136.140 32.060 139.770 33.260 ;
        RECT 136.140 31.010 137.640 32.060 ;
        RECT 137.900 31.700 138.130 32.060 ;
        RECT 138.340 31.650 139.390 31.710 ;
        RECT 139.540 31.700 139.770 32.060 ;
        RECT 138.335 31.420 139.390 31.650 ;
        RECT 138.340 31.410 139.390 31.420 ;
        RECT 137.900 31.010 138.130 31.370 ;
        RECT 139.540 31.010 139.770 31.370 ;
        RECT 139.940 31.060 142.240 43.560 ;
        RECT 142.890 43.110 143.940 43.410 ;
        RECT 136.140 29.810 139.770 31.010 ;
        RECT 136.140 29.160 137.640 29.810 ;
        RECT 137.900 29.410 138.130 29.810 ;
        RECT 139.540 29.410 139.770 29.810 ;
        RECT 138.615 29.360 139.165 29.390 ;
        RECT 131.940 29.110 137.640 29.160 ;
        RECT 126.950 27.940 127.180 28.360 ;
        RECT 127.340 27.610 128.340 27.960 ;
        RECT 126.950 27.210 127.180 27.610 ;
        RECT 128.490 27.210 129.440 28.360 ;
        RECT 133.140 28.210 137.640 29.110 ;
        RECT 138.290 29.060 139.390 29.360 ;
        RECT 138.390 28.810 139.340 29.060 ;
        RECT 138.615 28.780 139.165 28.810 ;
        RECT 133.140 27.410 135.490 28.210 ;
        RECT 138.340 27.710 139.340 28.110 ;
        RECT 132.240 27.300 135.490 27.410 ;
        RECT 136.790 27.460 139.340 27.710 ;
        RECT 136.790 27.300 139.190 27.460 ;
        RECT 140.390 27.410 142.240 31.060 ;
        RECT 142.390 30.310 142.740 43.110 ;
        RECT 144.140 42.620 144.370 43.080 ;
        RECT 142.940 42.570 143.990 42.610 ;
        RECT 142.935 42.340 143.990 42.570 ;
        RECT 142.940 42.310 143.990 42.340 ;
        RECT 144.740 42.510 149.340 42.660 ;
        RECT 150.790 42.510 153.090 92.010 ;
        RECT 144.740 42.500 153.350 42.510 ;
        RECT 144.140 41.830 144.370 42.290 ;
        RECT 142.890 41.510 143.940 41.810 ;
        RECT 144.740 41.700 155.700 42.500 ;
        RECT 144.140 41.040 144.370 41.500 ;
        RECT 142.940 40.990 143.990 41.010 ;
        RECT 142.935 40.760 143.990 40.990 ;
        RECT 142.940 40.710 143.990 40.760 ;
        RECT 144.740 40.800 157.310 41.700 ;
        RECT 142.890 39.960 143.940 40.260 ;
        RECT 144.140 40.250 144.370 40.710 ;
        RECT 144.740 40.210 155.700 40.800 ;
        RECT 156.410 40.600 157.310 40.800 ;
        RECT 144.140 39.460 144.370 39.920 ;
        RECT 144.740 39.460 149.340 40.210 ;
        RECT 152.660 40.200 155.700 40.210 ;
        RECT 156.380 39.700 157.340 40.600 ;
        RECT 142.940 39.410 143.990 39.460 ;
        RECT 142.935 39.180 143.990 39.410 ;
        RECT 142.940 39.160 143.990 39.180 ;
        RECT 144.740 39.410 148.090 39.460 ;
        RECT 144.140 38.670 144.370 39.130 ;
        RECT 142.890 38.360 143.940 38.660 ;
        RECT 144.140 37.880 144.370 38.340 ;
        RECT 142.940 37.830 143.990 37.860 ;
        RECT 142.935 37.600 143.990 37.830 ;
        RECT 142.940 37.560 143.990 37.600 ;
        RECT 144.140 37.090 144.370 37.550 ;
        RECT 142.890 36.760 143.940 37.060 ;
        RECT 144.140 36.300 144.370 36.760 ;
        RECT 142.940 36.250 143.990 36.260 ;
        RECT 142.935 36.020 143.990 36.250 ;
        RECT 142.940 35.960 143.990 36.020 ;
        RECT 144.140 35.510 144.370 35.970 ;
        RECT 142.890 35.210 143.940 35.510 ;
        RECT 144.140 34.720 144.370 35.180 ;
        RECT 142.940 34.670 143.990 34.710 ;
        RECT 142.935 34.440 143.990 34.670 ;
        RECT 142.940 34.410 143.990 34.440 ;
        RECT 144.140 33.930 144.370 34.390 ;
        RECT 142.890 33.610 143.940 33.910 ;
        RECT 142.940 33.090 143.990 33.160 ;
        RECT 144.140 33.140 144.370 33.600 ;
        RECT 142.935 32.860 143.990 33.090 ;
        RECT 142.890 32.060 143.940 32.360 ;
        RECT 144.140 32.350 144.370 32.810 ;
        RECT 144.140 31.560 144.370 32.020 ;
        RECT 142.940 31.510 143.990 31.560 ;
        RECT 142.935 31.280 143.990 31.510 ;
        RECT 142.940 31.260 143.990 31.280 ;
        RECT 144.140 30.770 144.370 31.230 ;
        RECT 142.890 30.460 143.940 30.760 ;
        RECT 142.390 29.410 142.790 30.310 ;
        RECT 144.140 29.980 144.370 30.440 ;
        RECT 142.940 29.930 143.990 29.960 ;
        RECT 142.935 29.700 143.990 29.930 ;
        RECT 142.940 29.660 143.990 29.700 ;
        RECT 142.390 27.560 142.740 29.410 ;
        RECT 144.140 29.190 144.370 29.650 ;
        RECT 142.890 28.860 143.940 29.160 ;
        RECT 142.940 28.350 143.990 28.410 ;
        RECT 144.140 28.400 144.370 28.860 ;
        RECT 142.935 28.120 143.990 28.350 ;
        RECT 142.940 28.110 143.990 28.120 ;
        RECT 144.140 27.610 144.370 28.070 ;
        RECT 142.890 27.310 143.940 27.610 ;
        RECT 126.940 26.060 129.440 27.210 ;
        RECT 130.240 26.870 131.240 27.260 ;
        RECT 132.090 27.160 135.490 27.300 ;
        RECT 132.090 27.070 134.590 27.160 ;
        RECT 136.690 27.070 139.190 27.300 ;
        RECT 132.240 27.060 134.540 27.070 ;
        RECT 131.700 26.960 131.930 27.020 ;
        RECT 134.750 26.960 134.980 27.020 ;
        RECT 136.300 26.960 136.530 27.020 ;
        RECT 139.350 26.960 139.580 27.020 ;
        RECT 131.590 26.870 131.990 26.960 ;
        RECT 134.690 26.870 135.090 26.960 ;
        RECT 130.240 26.655 135.090 26.870 ;
        RECT 130.240 26.260 131.240 26.655 ;
        RECT 131.590 26.610 131.990 26.655 ;
        RECT 134.690 26.610 135.090 26.655 ;
        RECT 136.190 26.885 136.590 26.960 ;
        RECT 139.290 26.885 139.690 26.960 ;
        RECT 140.090 26.885 141.090 27.260 ;
        RECT 136.190 26.660 141.090 26.885 ;
        RECT 136.190 26.610 136.590 26.660 ;
        RECT 139.290 26.640 141.090 26.660 ;
        RECT 139.290 26.610 139.690 26.640 ;
        RECT 131.700 26.560 131.930 26.610 ;
        RECT 134.750 26.560 134.980 26.610 ;
        RECT 136.300 26.560 136.530 26.610 ;
        RECT 139.350 26.560 139.580 26.610 ;
        RECT 132.090 26.410 134.590 26.510 ;
        RECT 136.690 26.410 139.190 26.510 ;
        RECT 132.090 26.280 139.190 26.410 ;
        RECT 132.290 26.060 138.940 26.280 ;
        RECT 140.090 26.260 141.090 26.640 ;
        RECT 144.740 26.610 146.040 39.410 ;
        RECT 146.840 39.260 147.890 39.410 ;
        RECT 146.890 39.160 147.890 39.260 ;
        RECT 146.500 38.760 146.730 39.110 ;
        RECT 146.390 38.560 146.740 38.760 ;
        RECT 148.050 38.560 148.280 39.110 ;
        RECT 146.390 37.610 148.280 38.560 ;
        RECT 146.390 36.310 146.740 37.610 ;
        RECT 146.890 36.860 147.890 37.160 ;
        RECT 148.050 37.150 148.280 37.610 ;
        RECT 148.050 36.310 148.280 36.820 ;
        RECT 146.390 35.360 148.280 36.310 ;
        RECT 146.390 33.960 146.740 35.360 ;
        RECT 148.050 34.860 148.280 35.360 ;
        RECT 146.890 34.560 147.890 34.860 ;
        RECT 148.050 33.960 148.280 34.530 ;
        RECT 146.390 33.010 148.280 33.960 ;
        RECT 146.390 31.810 146.740 33.010 ;
        RECT 148.050 32.570 148.280 33.010 ;
        RECT 146.890 32.260 147.890 32.560 ;
        RECT 148.050 31.810 148.280 32.240 ;
        RECT 146.390 30.860 148.280 31.810 ;
        RECT 146.390 29.510 146.740 30.860 ;
        RECT 146.890 29.960 147.890 30.310 ;
        RECT 148.050 30.280 148.280 30.860 ;
        RECT 148.050 29.510 148.280 29.950 ;
        RECT 146.390 28.560 148.280 29.510 ;
        RECT 146.390 27.260 146.740 28.560 ;
        RECT 146.890 27.660 147.890 28.010 ;
        RECT 148.050 27.990 148.280 28.560 ;
        RECT 148.050 27.260 148.280 27.660 ;
        RECT 146.390 26.310 148.280 27.260 ;
        RECT 126.950 25.650 127.180 26.060 ;
        RECT 128.490 25.810 129.440 26.060 ;
        RECT 128.490 25.660 129.820 25.810 ;
        RECT 131.140 25.660 132.140 25.960 ;
        RECT 127.340 25.360 129.820 25.660 ;
        RECT 126.950 24.960 127.180 25.320 ;
        RECT 128.490 25.160 129.820 25.360 ;
        RECT 128.490 24.960 129.440 25.160 ;
        RECT 133.140 25.110 138.390 26.060 ;
        RECT 139.290 25.660 140.290 25.960 ;
        RECT 144.245 25.930 145.135 25.960 ;
        RECT 146.390 25.930 146.740 26.310 ;
        RECT 144.245 25.040 146.740 25.930 ;
        RECT 148.050 25.700 148.280 26.310 ;
        RECT 146.990 25.650 147.890 25.660 ;
        RECT 146.890 25.420 147.890 25.650 ;
        RECT 146.990 25.360 147.890 25.420 ;
        RECT 144.245 25.010 145.135 25.040 ;
        RECT 126.940 23.810 129.440 24.960 ;
        RECT 146.390 24.910 146.740 25.040 ;
        RECT 148.050 24.910 148.280 25.370 ;
        RECT 131.340 24.620 133.300 24.850 ;
        RECT 133.630 24.620 135.590 24.850 ;
        RECT 135.920 24.620 137.880 24.850 ;
        RECT 138.210 24.620 140.170 24.850 ;
        RECT 131.060 24.410 131.290 24.460 ;
        RECT 126.950 23.360 127.180 23.810 ;
        RECT 128.490 23.360 129.440 23.810 ;
        RECT 130.940 23.510 131.340 24.410 ;
        RECT 131.060 23.460 131.290 23.510 ;
        RECT 128.540 23.310 129.440 23.360 ;
        RECT 131.790 23.310 132.690 24.620 ;
        RECT 133.350 24.310 133.580 24.460 ;
        RECT 133.240 23.610 133.690 24.310 ;
        RECT 133.350 23.460 133.580 23.610 ;
        RECT 134.190 23.310 135.090 24.620 ;
        RECT 135.640 24.310 135.870 24.460 ;
        RECT 135.540 23.610 135.990 24.310 ;
        RECT 135.640 23.460 135.870 23.610 ;
        RECT 136.490 23.310 137.390 24.620 ;
        RECT 137.930 24.310 138.160 24.460 ;
        RECT 137.840 23.610 138.290 24.310 ;
        RECT 137.930 23.460 138.160 23.610 ;
        RECT 138.740 23.310 139.640 24.620 ;
        RECT 140.220 24.410 140.450 24.460 ;
        RECT 140.140 23.510 140.540 24.410 ;
        RECT 140.220 23.460 140.450 23.510 ;
        RECT 127.340 22.960 128.340 23.310 ;
        RECT 128.540 23.300 140.140 23.310 ;
        RECT 128.540 23.070 140.170 23.300 ;
        RECT 128.540 23.010 140.140 23.070 ;
        RECT 140.740 22.810 142.090 24.860 ;
        RECT 144.540 22.810 146.240 24.310 ;
        RECT 146.390 23.960 148.340 24.910 ;
        RECT 148.590 24.310 149.340 37.260 ;
        RECT 146.390 23.460 146.740 23.960 ;
        RECT 146.500 23.410 146.730 23.460 ;
        RECT 148.050 23.410 148.280 23.960 ;
        RECT 146.890 23.060 147.890 23.410 ;
        RECT 148.490 22.810 149.340 24.310 ;
        RECT 125.140 21.605 149.340 22.810 ;
        RECT 105.470 20.460 149.340 21.605 ;
        RECT 105.470 20.415 118.640 20.460 ;
        RECT 122.640 20.415 130.285 20.460 ;
        RECT 115.540 20.410 116.290 20.415 ;
        RECT 115.770 18.310 116.020 18.625 ;
        RECT 119.820 18.310 120.070 18.825 ;
        RECT 115.540 17.110 120.340 18.310 ;
        RECT 115.770 16.520 116.020 17.110 ;
        RECT 117.340 14.860 118.540 17.110 ;
        RECT 119.820 16.720 120.070 17.110 ;
        RECT 150.940 14.860 152.140 14.890 ;
        RECT 117.340 13.660 152.140 14.860 ;
        RECT 150.940 13.630 152.140 13.660 ;
      LAYER via ;
        RECT 102.780 90.345 103.805 91.370 ;
        RECT 127.110 88.700 127.790 89.380 ;
        RECT 111.765 68.055 112.955 69.245 ;
        RECT 147.090 82.020 148.190 83.120 ;
        RECT 112.490 67.010 113.210 67.730 ;
        RECT 144.780 48.580 145.700 49.500 ;
        RECT 138.340 42.860 139.340 43.160 ;
        RECT 129.890 40.860 130.740 41.210 ;
        RECT 129.790 40.560 130.740 40.860 ;
        RECT 125.290 22.910 126.090 32.710 ;
        RECT 127.390 32.210 128.290 32.560 ;
        RECT 129.890 36.260 130.740 40.560 ;
        RECT 129.790 35.960 130.740 36.260 ;
        RECT 129.890 31.710 130.740 35.960 ;
        RECT 129.790 31.410 130.740 31.710 ;
        RECT 129.890 31.260 130.740 31.410 ;
        RECT 132.040 40.560 132.940 40.860 ;
        RECT 132.040 35.960 132.940 36.260 ;
        RECT 132.040 31.410 132.940 31.710 ;
        RECT 138.440 40.560 139.340 40.860 ;
        RECT 138.340 38.260 139.340 38.560 ;
        RECT 138.440 35.960 139.340 36.260 ;
        RECT 138.340 33.660 139.340 33.960 ;
        RECT 138.440 31.410 139.340 31.710 ;
        RECT 140.640 33.960 141.490 43.610 ;
        RECT 142.940 43.110 143.890 43.410 ;
        RECT 140.640 33.560 141.540 33.960 ;
        RECT 140.640 32.410 141.490 33.560 ;
        RECT 140.640 32.010 141.540 32.410 ;
        RECT 127.390 27.610 128.290 27.960 ;
        RECT 138.340 29.060 139.340 29.360 ;
        RECT 138.615 28.810 139.165 29.060 ;
        RECT 138.390 27.460 139.240 28.110 ;
        RECT 140.640 30.810 141.490 32.010 ;
        RECT 140.640 27.810 141.540 30.810 ;
        RECT 140.640 27.460 141.890 27.810 ;
        RECT 140.740 27.410 141.890 27.460 ;
        RECT 142.990 42.310 143.940 42.610 ;
        RECT 142.940 41.510 143.890 41.810 ;
        RECT 142.990 40.710 143.940 41.010 ;
        RECT 142.940 39.960 143.890 40.260 ;
        RECT 142.990 39.160 143.940 39.460 ;
        RECT 142.940 38.360 143.890 38.660 ;
        RECT 142.990 37.560 143.940 37.860 ;
        RECT 142.940 36.760 143.890 37.060 ;
        RECT 142.990 35.960 143.940 36.260 ;
        RECT 142.940 35.210 143.890 35.510 ;
        RECT 142.990 34.410 143.940 34.710 ;
        RECT 142.940 33.610 143.890 33.910 ;
        RECT 142.990 32.860 143.940 33.160 ;
        RECT 142.940 32.060 143.890 32.360 ;
        RECT 142.990 31.260 143.940 31.560 ;
        RECT 142.940 30.460 143.890 30.760 ;
        RECT 142.440 29.610 142.740 30.010 ;
        RECT 142.990 29.660 143.940 29.960 ;
        RECT 142.940 28.860 143.890 29.160 ;
        RECT 142.990 28.110 143.940 28.410 ;
        RECT 142.940 27.310 143.890 27.610 ;
        RECT 130.340 27.040 131.040 27.060 ;
        RECT 130.315 26.485 131.040 27.040 ;
        RECT 130.340 26.460 131.040 26.485 ;
        RECT 131.640 26.610 131.940 26.960 ;
        RECT 134.740 26.610 135.040 26.960 ;
        RECT 136.240 26.610 136.540 26.960 ;
        RECT 139.340 26.610 139.640 26.960 ;
        RECT 140.365 26.490 140.915 27.040 ;
        RECT 145.090 26.610 145.690 42.460 ;
        RECT 148.790 39.760 149.190 42.460 ;
        RECT 156.410 39.700 157.310 40.600 ;
        RECT 146.890 39.260 147.840 39.560 ;
        RECT 147.040 39.160 147.790 39.260 ;
        RECT 146.940 36.860 147.840 37.160 ;
        RECT 146.940 34.560 147.840 34.860 ;
        RECT 146.940 32.260 147.840 32.560 ;
        RECT 146.940 29.960 147.840 30.310 ;
        RECT 146.940 27.660 147.840 28.010 ;
        RECT 129.140 25.160 129.790 25.810 ;
        RECT 131.190 25.660 132.090 25.960 ;
        RECT 133.290 25.410 133.690 26.110 ;
        RECT 137.840 25.410 138.240 26.110 ;
        RECT 139.340 25.660 140.240 25.960 ;
        RECT 147.040 25.360 147.840 25.660 ;
        RECT 130.990 23.510 131.290 24.410 ;
        RECT 133.290 23.610 133.640 24.310 ;
        RECT 135.590 23.610 135.940 24.310 ;
        RECT 137.890 23.610 138.240 24.310 ;
        RECT 140.190 23.510 140.490 24.410 ;
        RECT 127.390 22.960 128.290 23.310 ;
        RECT 148.740 24.610 149.140 37.110 ;
        RECT 146.940 23.060 147.840 23.410 ;
        RECT 130.840 22.260 131.340 22.360 ;
        RECT 135.590 22.260 135.940 22.360 ;
        RECT 139.990 22.260 140.490 22.360 ;
        RECT 130.840 21.910 140.490 22.260 ;
        RECT 130.840 21.610 140.440 21.910 ;
        RECT 150.940 13.660 152.140 14.860 ;
      LAYER met2 ;
        RECT 102.780 89.445 103.805 91.400 ;
        RECT 102.760 88.470 103.825 89.445 ;
        RECT 102.780 88.445 103.805 88.470 ;
        RECT 127.110 87.575 127.790 89.410 ;
        RECT 90.275 83.250 91.725 83.270 ;
        RECT 90.250 81.750 95.280 83.250 ;
        RECT 90.275 81.730 91.725 81.750 ;
        RECT 147.090 79.605 148.190 83.150 ;
        RECT 147.070 78.555 148.210 79.605 ;
        RECT 147.090 78.530 148.190 78.555 ;
        RECT 111.765 69.245 112.955 69.275 ;
        RECT 111.765 68.055 114.840 69.245 ;
        RECT 111.765 68.025 112.955 68.055 ;
        RECT 107.760 67.730 108.480 67.775 ;
        RECT 112.490 67.730 113.210 67.760 ;
        RECT 107.760 67.010 113.210 67.730 ;
        RECT 107.760 66.965 108.480 67.010 ;
        RECT 112.490 66.980 113.210 67.010 ;
        RECT 144.750 49.475 146.470 49.500 ;
        RECT 144.750 48.605 146.490 49.475 ;
        RECT 144.750 48.580 146.470 48.605 ;
        RECT 66.775 45.250 68.225 45.270 ;
        RECT 98.970 45.250 112.970 45.260 ;
        RECT 66.750 43.760 112.970 45.250 ;
        RECT 66.750 43.750 99.710 43.760 ;
        RECT 66.775 43.730 68.225 43.750 ;
        RECT 140.640 43.460 141.490 43.660 ;
        RECT 134.750 43.410 136.530 43.450 ;
        RECT 134.740 43.160 139.390 43.410 ;
        RECT 134.750 42.860 139.390 43.160 ;
        RECT 140.640 43.060 143.940 43.460 ;
        RECT 134.750 42.820 139.340 42.860 ;
        RECT 129.890 40.910 130.740 41.260 ;
        RECT 129.790 40.860 130.740 40.910 ;
        RECT 132.040 40.860 132.940 40.910 ;
        RECT 129.740 40.560 133.190 40.860 ;
        RECT 129.790 40.510 130.740 40.560 ;
        RECT 132.040 40.510 132.940 40.560 ;
        RECT 129.890 36.310 130.740 40.510 ;
        RECT 134.750 38.600 136.530 42.820 ;
        RECT 138.340 42.810 139.340 42.820 ;
        RECT 140.640 41.860 141.490 43.060 ;
        RECT 142.940 42.260 149.340 42.660 ;
        RECT 140.640 41.460 143.940 41.860 ;
        RECT 140.640 40.910 141.490 41.460 ;
        RECT 144.740 41.010 149.340 42.260 ;
        RECT 138.440 40.560 141.490 40.910 ;
        RECT 142.940 40.710 149.340 41.010 ;
        RECT 138.440 40.510 139.340 40.560 ;
        RECT 140.640 40.310 141.490 40.560 ;
        RECT 140.640 39.910 143.940 40.310 ;
        RECT 140.640 38.710 141.490 39.910 ;
        RECT 144.790 39.460 149.340 40.710 ;
        RECT 142.940 39.160 148.040 39.460 ;
        RECT 144.740 39.010 148.040 39.160 ;
        RECT 138.340 38.600 139.340 38.610 ;
        RECT 134.750 38.220 139.390 38.600 ;
        RECT 140.640 38.310 143.940 38.710 ;
        RECT 129.790 36.260 130.740 36.310 ;
        RECT 132.040 36.260 132.940 36.310 ;
        RECT 129.740 35.960 133.190 36.260 ;
        RECT 129.790 35.910 130.740 35.960 ;
        RECT 132.040 35.910 132.940 35.960 ;
        RECT 125.290 32.710 126.090 32.760 ;
        RECT 125.290 32.060 128.440 32.710 ;
        RECT 125.290 28.160 126.090 32.060 ;
        RECT 129.890 31.760 130.740 35.910 ;
        RECT 134.750 34.000 136.530 38.220 ;
        RECT 138.340 38.210 139.340 38.220 ;
        RECT 140.640 37.110 141.490 38.310 ;
        RECT 144.740 37.860 146.040 39.010 ;
        RECT 142.940 37.560 146.040 37.860 ;
        RECT 140.640 36.710 143.890 37.110 ;
        RECT 140.640 36.360 141.490 36.710 ;
        RECT 138.440 35.960 141.490 36.360 ;
        RECT 144.740 36.310 146.040 37.560 ;
        RECT 146.890 36.710 149.340 37.260 ;
        RECT 142.940 35.960 146.040 36.310 ;
        RECT 138.440 35.910 139.340 35.960 ;
        RECT 140.640 35.560 141.490 35.960 ;
        RECT 140.640 35.160 143.890 35.560 ;
        RECT 138.340 34.000 139.340 34.010 ;
        RECT 134.750 33.620 139.340 34.000 ;
        RECT 129.790 31.710 130.740 31.760 ;
        RECT 132.040 31.710 132.940 31.760 ;
        RECT 129.740 31.410 133.190 31.710 ;
        RECT 129.790 31.360 130.740 31.410 ;
        RECT 132.040 31.360 132.940 31.410 ;
        RECT 129.890 31.210 130.740 31.360 ;
        RECT 134.750 30.120 136.530 33.620 ;
        RECT 138.340 33.610 139.340 33.620 ;
        RECT 140.640 33.960 141.490 35.160 ;
        RECT 144.740 34.960 146.040 35.960 ;
        RECT 144.740 34.710 148.040 34.960 ;
        RECT 142.940 34.410 148.040 34.710 ;
        RECT 142.940 34.360 146.040 34.410 ;
        RECT 140.640 33.560 143.940 33.960 ;
        RECT 140.640 32.410 141.490 33.560 ;
        RECT 144.740 33.160 146.040 34.360 ;
        RECT 142.940 32.810 146.040 33.160 ;
        RECT 140.640 32.010 143.940 32.410 ;
        RECT 140.640 31.760 141.490 32.010 ;
        RECT 138.440 31.410 141.490 31.760 ;
        RECT 144.740 31.560 146.040 32.810 ;
        RECT 148.590 32.710 149.340 36.710 ;
        RECT 156.410 34.925 157.310 40.630 ;
        RECT 156.390 34.075 157.330 34.925 ;
        RECT 156.410 34.050 157.310 34.075 ;
        RECT 146.890 32.160 149.340 32.710 ;
        RECT 138.440 31.360 139.340 31.410 ;
        RECT 140.640 30.810 141.490 31.410 ;
        RECT 142.940 31.210 146.040 31.560 ;
        RECT 140.640 30.410 143.940 30.810 ;
        RECT 134.760 28.880 136.520 30.120 ;
        RECT 138.615 29.410 139.165 29.980 ;
        RECT 125.290 27.510 128.440 28.160 ;
        RECT 138.340 27.860 139.340 29.410 ;
        RECT 140.640 29.210 141.540 30.410 ;
        RECT 144.740 30.360 146.040 31.210 ;
        RECT 141.740 29.560 142.740 30.060 ;
        RECT 144.740 30.010 148.040 30.360 ;
        RECT 142.940 29.810 148.040 30.010 ;
        RECT 142.940 29.610 146.040 29.810 ;
        RECT 141.740 29.510 142.440 29.560 ;
        RECT 140.640 28.810 143.890 29.210 ;
        RECT 140.640 27.860 141.540 28.810 ;
        RECT 144.740 28.460 146.040 29.610 ;
        RECT 142.940 28.060 146.040 28.460 ;
        RECT 148.590 28.110 149.340 32.160 ;
        RECT 125.290 23.560 126.090 27.510 ;
        RECT 129.940 27.040 131.140 27.760 ;
        RECT 138.390 27.410 139.240 27.860 ;
        RECT 140.640 27.710 141.890 27.860 ;
        RECT 140.640 27.410 143.890 27.710 ;
        RECT 141.790 27.260 143.890 27.410 ;
        RECT 140.290 27.040 141.590 27.260 ;
        RECT 129.940 27.010 135.015 27.040 ;
        RECT 136.265 27.010 141.590 27.040 ;
        RECT 129.940 26.560 135.040 27.010 ;
        RECT 136.240 26.560 141.590 27.010 ;
        RECT 144.740 27.210 146.040 28.060 ;
        RECT 146.890 27.560 149.340 28.110 ;
        RECT 144.740 26.610 147.840 27.210 ;
        RECT 129.940 26.485 135.015 26.560 ;
        RECT 136.265 26.490 141.590 26.560 ;
        RECT 129.940 26.310 131.140 26.485 ;
        RECT 140.290 26.260 141.590 26.490 ;
        RECT 129.140 25.810 129.790 25.840 ;
        RECT 129.140 25.160 130.510 25.810 ;
        RECT 130.790 25.560 132.140 26.010 ;
        RECT 129.140 25.130 129.790 25.160 ;
        RECT 125.290 22.910 128.440 23.560 ;
        RECT 125.290 22.860 126.090 22.910 ;
        RECT 130.790 22.360 131.440 25.560 ;
        RECT 133.190 23.460 133.790 26.210 ;
        RECT 135.490 22.360 136.040 24.460 ;
        RECT 137.740 23.460 138.340 26.210 ;
        RECT 139.240 25.560 140.590 26.010 ;
        RECT 143.225 25.930 144.065 26.105 ;
        RECT 139.940 22.360 140.590 25.560 ;
        RECT 143.200 25.040 145.165 25.930 ;
        RECT 147.040 25.310 147.840 26.610 ;
        RECT 143.225 24.865 144.065 25.040 ;
        RECT 148.590 23.560 149.340 27.560 ;
        RECT 146.890 23.010 149.340 23.560 ;
        RECT 130.790 21.460 140.590 22.360 ;
        RECT 150.940 14.860 152.140 22.155 ;
        RECT 150.910 13.660 152.170 14.860 ;
      LAYER via2 ;
        RECT 102.805 88.470 103.780 89.445 ;
        RECT 127.110 87.620 127.790 88.300 ;
        RECT 90.275 81.775 91.725 83.225 ;
        RECT 147.115 78.555 148.165 79.605 ;
        RECT 113.605 68.055 114.795 69.245 ;
        RECT 145.575 48.605 146.445 49.475 ;
        RECT 66.775 43.775 68.225 45.225 ;
        RECT 156.435 34.075 157.285 34.925 ;
        RECT 134.990 29.360 136.440 30.160 ;
        RECT 138.615 29.385 139.165 29.935 ;
        RECT 130.040 27.110 130.640 27.660 ;
        RECT 140.890 26.460 141.490 27.160 ;
        RECT 129.815 25.160 130.465 25.810 ;
        RECT 143.225 24.910 144.065 26.060 ;
        RECT 150.940 20.910 152.140 22.110 ;
      LAYER met3 ;
        RECT 87.255 83.250 88.745 83.275 ;
        RECT 87.250 81.750 91.750 83.250 ;
        RECT 87.255 81.725 88.745 81.750 ;
        RECT 28.255 45.250 29.745 45.275 ;
        RECT 28.250 43.750 68.250 45.250 ;
        RECT 28.255 43.725 29.745 43.750 ;
        RECT 102.780 27.510 103.805 89.470 ;
        RECT 127.085 87.595 127.815 88.325 ;
        RECT 127.110 86.800 127.790 87.595 ;
        RECT 110.070 70.460 126.930 85.860 ;
        RECT 128.770 69.750 145.630 85.150 ;
        RECT 113.580 69.245 114.820 69.270 ;
        RECT 113.580 68.055 116.365 69.245 ;
        RECT 113.580 68.030 114.820 68.055 ;
        RECT 147.090 67.995 148.190 79.630 ;
        RECT 107.735 66.985 108.505 67.755 ;
        RECT 107.760 63.150 108.480 66.985 ;
        RECT 109.980 51.340 126.840 66.740 ;
        RECT 128.940 51.540 145.800 66.940 ;
        RECT 147.065 66.905 148.215 67.995 ;
        RECT 147.090 66.900 148.190 66.905 ;
        RECT 145.550 50.065 146.470 50.070 ;
        RECT 145.525 49.155 146.495 50.065 ;
        RECT 145.550 48.580 146.470 49.155 ;
        RECT 134.890 30.175 141.840 30.210 ;
        RECT 134.890 29.985 142.405 30.175 ;
        RECT 134.890 29.535 142.440 29.985 ;
        RECT 134.890 29.350 142.405 29.535 ;
        RECT 134.890 29.260 141.840 29.350 ;
        RECT 137.190 28.760 140.040 29.260 ;
        RECT 123.990 27.510 130.840 27.860 ;
        RECT 102.780 26.960 130.840 27.510 ;
        RECT 140.840 27.310 150.690 27.410 ;
        RECT 102.780 26.510 124.640 26.960 ;
        RECT 140.840 26.610 152.140 27.310 ;
        RECT 102.780 26.500 103.805 26.510 ;
        RECT 140.840 26.410 141.640 26.610 ;
        RECT 149.840 26.110 152.140 26.610 ;
        RECT 129.540 24.885 144.090 26.085 ;
        RECT 150.940 22.135 152.140 26.110 ;
        RECT 150.915 20.885 152.165 22.135 ;
        RECT 156.410 8.645 157.310 34.950 ;
        RECT 156.385 7.755 157.335 8.645 ;
        RECT 156.410 7.750 157.310 7.755 ;
      LAYER via3 ;
        RECT 87.255 81.755 88.745 83.245 ;
        RECT 28.255 43.755 29.745 45.245 ;
        RECT 127.110 86.830 127.790 87.510 ;
        RECT 126.510 70.600 126.830 85.720 ;
        RECT 145.210 69.890 145.530 85.010 ;
        RECT 115.145 68.055 116.335 69.245 ;
        RECT 147.095 66.905 148.185 67.995 ;
        RECT 107.760 63.180 108.480 63.900 ;
        RECT 126.420 51.480 126.740 66.600 ;
        RECT 145.380 51.680 145.700 66.800 ;
        RECT 145.555 49.155 146.465 50.065 ;
        RECT 156.415 7.755 157.305 8.645 ;
      LAYER met4 ;
        RECT 3.990 223.800 4.290 224.760 ;
        RECT 7.670 223.800 7.970 224.760 ;
        RECT 11.350 223.800 11.650 224.760 ;
        RECT 15.030 223.800 15.330 224.760 ;
        RECT 18.710 223.800 19.010 224.760 ;
        RECT 22.390 223.800 22.690 224.760 ;
        RECT 26.070 223.800 26.370 224.760 ;
        RECT 29.750 223.800 30.050 224.760 ;
        RECT 33.430 223.800 33.730 224.760 ;
        RECT 37.110 223.800 37.410 224.760 ;
        RECT 40.790 223.800 41.090 224.760 ;
        RECT 44.470 223.800 44.770 224.760 ;
        RECT 48.150 223.800 48.450 224.760 ;
        RECT 51.830 223.800 52.130 224.760 ;
        RECT 55.510 223.800 55.810 224.760 ;
        RECT 59.190 223.800 59.490 224.760 ;
        RECT 62.870 223.800 63.170 224.760 ;
        RECT 66.550 223.800 66.850 224.760 ;
        RECT 70.230 223.800 70.530 224.760 ;
        RECT 73.910 223.800 74.210 224.760 ;
        RECT 77.590 223.800 77.890 224.760 ;
        RECT 81.270 223.800 81.570 224.760 ;
        RECT 84.950 223.800 85.250 224.760 ;
        RECT 88.630 223.800 88.930 224.760 ;
        RECT 3.200 223.500 88.930 223.800 ;
        RECT 49.000 220.760 50.500 223.500 ;
        RECT 66.550 223.450 66.850 223.500 ;
        RECT 84.950 223.450 85.250 223.500 ;
        RECT 127.105 87.020 127.795 87.515 ;
        RECT 125.990 85.840 145.960 87.020 ;
        RECT 50.500 81.750 88.750 83.250 ;
        RECT 110.465 70.855 125.075 85.465 ;
        RECT 125.990 80.000 127.170 85.840 ;
        RECT 116.860 69.285 117.990 70.855 ;
        RECT 126.430 70.520 126.910 80.000 ;
        RECT 129.165 70.145 143.775 84.755 ;
        RECT 144.780 79.440 145.960 85.840 ;
        RECT 136.855 69.285 137.985 70.145 ;
        RECT 145.130 69.810 145.610 79.440 ;
        RECT 115.140 69.245 116.340 69.250 ;
        RECT 116.860 69.245 137.985 69.285 ;
        RECT 115.140 68.155 137.985 69.245 ;
        RECT 115.140 68.055 117.785 68.155 ;
        RECT 115.140 68.050 116.340 68.055 ;
        RECT 144.950 66.900 148.190 68.000 ;
        RECT 107.755 63.900 108.485 63.905 ;
        RECT 110.375 63.900 124.985 66.345 ;
        RECT 126.340 66.220 126.820 66.680 ;
        RECT 129.335 66.220 143.945 66.545 ;
        RECT 107.755 63.180 124.985 63.900 ;
        RECT 107.755 63.175 108.485 63.180 ;
        RECT 110.375 51.735 124.985 63.180 ;
        RECT 126.100 61.410 143.945 66.220 ;
        RECT 144.950 62.060 146.050 66.900 ;
        RECT 126.340 51.400 126.820 61.410 ;
        RECT 127.380 50.790 128.300 61.410 ;
        RECT 129.335 51.935 143.945 61.410 ;
        RECT 145.300 51.600 145.780 62.060 ;
        RECT 127.380 49.870 146.470 50.790 ;
        RECT 145.550 49.150 146.470 49.870 ;
        RECT 2.500 43.750 29.750 45.250 ;
        RECT 156.410 1.000 157.310 8.650 ;
  END
END tt_um_twin_tee_opamp_osc
END LIBRARY

