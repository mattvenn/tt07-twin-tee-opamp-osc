* NGSPICE file created from twin_tee_osc_parax.ext - technology: sky130A

.subckt twin_tee_osc_parax vdd vss out
X0 a_24144_17782# out.t18 vss.t28 sky130_fd_pr__res_high_po_0p35 l=50.36
X1 vss.t5 p3_opamp_0.PLUS vss.t4 sky130_fd_pr__res_high_po_0p35 l=20.16
X2 twin_tee_0.in.t1 twin_tee_0.c3_c4.t0 sky130_fd_pr__cap_mim_m3_1 l=15 w=15
X3 p3_opamp_0.VX p3_opamp_0.VBIAS.t9 vss.t8 vss.t7 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X4 vdd.t58 p3_opamp_0.V1.t7 out.t0 vdd.t57 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 vss.t12 twin_tee_0.c3_c4.t1 vss.t11 sky130_fd_pr__res_high_po_0p35 l=23.16
X6 vss.t10 p3_opamp_0.VBIAS.t10 p3_opamp_0.VX vss.t9 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X7 p3_opamp_0.VBIAS.t8 p3_opamp_0.VBIAS.t7 vss.t1 vss.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=2
X8 vss.t27 p3_opamp_0.VBIAS.t5 p3_opamp_0.VBIAS.t6 vss.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X9 vdd.t18 p3_opamp_0.VBIAS.t0 vss.t6 sky130_fd_pr__res_xhigh_po_0p35 l=2.88
X10 vdd.t56 p3_opamp_0.V1.t8 out.t23 vdd.t55 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X11 vdd.t9 p3_opamp_0.V2.t11 p3_opamp_0.V2.t12 vdd.t8 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=2
X12 p3_opamp_0.V2.t10 p3_opamp_0.V2.t9 vdd.t15 vdd.t14 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X13 twin_tee_0.in.t0 a_24144_17782# vss.t36 sky130_fd_pr__res_high_po_0p35 l=50.36
X14 vdd.t61 p3_opamp_0.V2.t7 p3_opamp_0.V2.t8 vdd.t60 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X15 vdd.t7 p3_opamp_0.V2.t13 p3_opamp_0.V1.t4 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=2
X16 out.t9 p3_opamp_0.V1.t9 vdd.t54 vdd.t53 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X17 p3_opamp_0.VX p3_opamp_0.VBIAS.t11 vss.t20 vss.t19 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=2
X18 vdd.t59 p3_opamp_0.PLUS vss.t18 sky130_fd_pr__res_high_po_0p35 l=20.16
X19 vdd.t3 p3_opamp_0.V2.t14 p3_opamp_0.V1.t2 vdd.t2 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X20 p3_opamp_0.V1.t1 p3_opamp_0.V2.t15 vdd.t1 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X21 vss.t26 p3_opamp_0.VBIAS.t12 p3_opamp_0.VX vss.t25 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=2
X22 out.t15 p3_opamp_0.VBIAS.t13 vss.t24 vss.t23 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=2
X23 p3_opamp_0.VBIAS.t4 p3_opamp_0.VBIAS.t3 vss.t2 vss.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X24 p3_opamp_0.V2.t0 twin_tee_0.in.t2 p3_opamp_0.VX vss.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=0.5
X25 vdd.t52 p3_opamp_0.V1.t10 out.t12 vdd.t51 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X26 twin_tee_0.c3_c4.t2 out.t1 sky130_fd_pr__cap_mim_m3_1 l=15 w=15
X27 vdd.t50 p3_opamp_0.V1.t11 out.t25 vdd.t49 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X28 out.t14 p3_opamp_0.VBIAS.t14 vss.t22 vss.t21 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X29 vss.t30 p3_opamp_0.VBIAS.t15 out.t19 vss.t29 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X30 vss.t33 p3_opamp_0.VBIAS.t1 p3_opamp_0.VBIAS.t2 vss.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=2
X31 out.t4 p3_opamp_0.V1.t12 vdd.t48 vdd.t47 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X32 vdd.t46 p3_opamp_0.V1.t13 out.t2 vdd.t45 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X33 out.t17 p3_opamp_0.V1.t14 vdd.t44 vdd.t43 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X34 vdd.t13 p3_opamp_0.V2.t5 p3_opamp_0.V2.t6 vdd.t12 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X35 vdd.t42 p3_opamp_0.V1.t15 out.t6 vdd.t41 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X36 out.t21 p3_opamp_0.V1.t16 vdd.t40 vdd.t39 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X37 p3_opamp_0.V2.t4 p3_opamp_0.V2.t3 vdd.t65 vdd.t64 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=2
X38 p3_opamp_0.V2.t2 p3_opamp_0.V2.t1 vdd.t17 vdd.t16 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X39 vdd.t38 p3_opamp_0.V1.t17 out.t5 vdd.t37 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X40 out.t24 p3_opamp_0.V1.t18 vdd.t36 vdd.t35 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X41 vdd.t5 p3_opamp_0.V2.t16 p3_opamp_0.V1.t3 vdd.t4 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X42 vdd.t34 p3_opamp_0.V1.t19 out.t3 vdd.t33 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X43 out.t11 p3_opamp_0.V1.t20 vdd.t32 vdd.t31 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X44 p3_opamp_0.V1.t6 p3_opamp_0.V2.t17 vdd.t63 vdd.t62 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X45 out.t10 p3_opamp_0.V1.t21 vdd.t30 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X46 p3_opamp_0.V1.t5 p3_opamp_0.V2.t18 vdd.t11 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=2
X47 vdd.t28 p3_opamp_0.V1.t22 out.t13 vdd.t27 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X48 out.t20 p3_opamp_0.V1.t23 vdd.t26 vdd.t25 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X49 vss.t32 p3_opamp_0.VBIAS.t16 out.t22 vss.t31 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X50 out.t27 p3_opamp_0.VBIAS.t17 vss.t35 vss.t34 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X51 p3_opamp_0.V1.t0 p3_opamp_0.PLUS p3_opamp_0.VX vss.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=0.5
X52 out.t28 p3_opamp_0.V1.t24 vdd.t24 vdd.t23 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X53 out.t8 p3_opamp_0.VBIAS.t18 vss.t16 vss.t15 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=2
X54 vss.t14 p3_opamp_0.VBIAS.t19 out.t7 vss.t13 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X55 vss.t37 a_24144_17782# sky130_fd_pr__cap_mim_m3_1 l=15 w=15
X56 out.t16 p3_opamp_0.V1.t25 vdd.t22 vdd.t21 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X57 vdd.t20 p3_opamp_0.V1.t26 out.t26 vdd.t19 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X58 vss.t38 a_24144_17782# sky130_fd_pr__cap_mim_m3_1 l=15 w=15
R0 out.n6 out.n5 203.756
R1 out.n6 out.n4 203.499
R2 out.n28 out.n8 201.875
R3 out.n27 out.n9 201.695
R4 out.n24 out.n12 201.619
R5 out.n22 out.n14 201.619
R6 out.n23 out.n13 201.619
R7 out.n26 out.n10 201.619
R8 out.n19 out.n17 201.561
R9 out.n20 out.n16 201.561
R10 out.n7 out.t8 83.7297
R11 out.n19 out.n18 69.1449
R12 out.n21 out.n15 68.1265
R13 out.n25 out.n11 68.1259
R14 out.n0 out.t18 44.2614
R15 out.n12 out.t25 28.5655
R16 out.n12 out.t16 28.5655
R17 out.n17 out.t26 28.5655
R18 out.n17 out.t11 28.5655
R19 out.n16 out.t0 28.5655
R20 out.n16 out.t28 28.5655
R21 out.n14 out.t6 28.5655
R22 out.n14 out.t24 28.5655
R23 out.n13 out.t3 28.5655
R24 out.n13 out.t20 28.5655
R25 out.n10 out.t5 28.5655
R26 out.n10 out.t10 28.5655
R27 out.n9 out.t13 28.5655
R28 out.n9 out.t17 28.5655
R29 out.n8 out.t2 28.5655
R30 out.n8 out.t9 28.5655
R31 out.n5 out.t12 28.5655
R32 out.n5 out.t4 28.5655
R33 out.n4 out.t23 28.5655
R34 out.n4 out.t21 28.5655
R35 out.n11 out.t22 17.4005
R36 out.n11 out.t14 17.4005
R37 out.n15 out.t7 17.4005
R38 out.n15 out.t27 17.4005
R39 out.n18 out.t19 17.4005
R40 out.n18 out.t15 17.4005
R41 out.n0 out.t1 4.93405
R42 out.n31 out.n2 2.69072
R43 out.n2 out 2.15883
R44 out.n29 out.n7 1.38826
R45 out.n30 out.n29 0.663586
R46 out.n24 out 0.565168
R47 out.n29 out.n28 0.285222
R48 out.n2 out.n1 0.17767
R49 out.n23 out.n22 0.154346
R50 out.n27 out.n26 0.151942
R51 out.n24 out.n23 0.149538
R52 out.n20 out.n19 0.149538
R53 out.n26 out.n25 0.139923
R54 out.n28 out.n27 0.1255
R55 out.n22 out.n21 0.1255
R56 out out.n31 0.1255
R57 out out.n30 0.0929762
R58 out.n1 out 0.0713874
R59 out.n29 out.n6 0.0639766
R60 out.n30 out.n3 0.0635409
R61 out.n31 out 0.063
R62 out.n1 out 0.0609244
R63 out.n21 out.n20 0.0269423
R64 out out.n3 0.0264615
R65 out out.n0 0.0167338
R66 out.n25 out.n24 0.0149231
R67 out.n7 out.n3 0.00499257
R68 vss.n65 vss.n64 258162
R69 vss.n64 vss.n63 140742
R70 vss.n66 vss.n65 92686.6
R71 vss.n64 vss.n32 21457
R72 vss.n155 vss.n149 17243.3
R73 vss.n155 vss.n150 17243.3
R74 vss.n149 vss.n6 17243.3
R75 vss.n150 vss.n6 17243.3
R76 vss.n78 vss.n44 15505.1
R77 vss.n74 vss.n44 15505.1
R78 vss.n78 vss.n45 15505.1
R79 vss.n74 vss.n45 15505.1
R80 vss.n71 vss.n47 15505.1
R81 vss.n67 vss.n47 15505.1
R82 vss.n71 vss.n48 15505.1
R83 vss.n67 vss.n48 15505.1
R84 vss.n137 vss.n7 11339.1
R85 vss.n50 vss.n7 11339.1
R86 vss.n137 vss.n8 11339.1
R87 vss.n50 vss.n8 11339.1
R88 vss.n146 vss.n139 9595.06
R89 vss.n142 vss.n139 9595.06
R90 vss.n146 vss.n140 9595.06
R91 vss.n142 vss.n140 9595.06
R92 vss.n157 vss.n2 9595.06
R93 vss.n161 vss.n2 9595.06
R94 vss.n157 vss.n3 9595.06
R95 vss.n161 vss.n3 9595.06
R96 vss.n122 vss.n29 7358.53
R97 vss.n122 vss.n30 7358.53
R98 vss.n124 vss.n30 7358.53
R99 vss.n124 vss.n29 7358.53
R100 vss.n81 vss.n35 7358.53
R101 vss.n81 vss.n36 7358.53
R102 vss.n117 vss.n36 7358.53
R103 vss.n117 vss.n35 7358.53
R104 vss.n114 vss.n38 5492.82
R105 vss.n114 vss.n39 5492.82
R106 vss.n42 vss.n38 5492.82
R107 vss.n42 vss.n39 5492.82
R108 vss.n90 vss.n87 3377.97
R109 vss.n93 vss.n87 3377.97
R110 vss.n90 vss.n88 3377.97
R111 vss.n93 vss.n88 3377.97
R112 vss.n60 vss.n52 3377.97
R113 vss.n55 vss.n52 3377.97
R114 vss.n60 vss.n53 3377.97
R115 vss.n55 vss.n53 3377.97
R116 vss.n148 vss.n138 2707.5
R117 vss.t31 vss.t15 1211.06
R118 vss.t21 vss.t31 1211.06
R119 vss.t13 vss.t21 1211.06
R120 vss.t34 vss.t13 1211.06
R121 vss.t29 vss.t34 1211.06
R122 vss.n63 vss.n51 1186.59
R123 vss.n154 vss.n151 1120.38
R124 vss.n154 vss.n153 1120.38
R125 vss.n152 vss.n151 1120.38
R126 vss.n153 vss.n152 1120.38
R127 vss.n77 vss.n46 1007.44
R128 vss.n75 vss.n46 1007.44
R129 vss.n77 vss.n76 1007.44
R130 vss.n76 vss.n75 1007.44
R131 vss.n70 vss.n49 1007.44
R132 vss.n68 vss.n49 1007.44
R133 vss.n70 vss.n69 1007.44
R134 vss.n69 vss.n68 1007.44
R135 vss.n138 vss.t15 906.971
R136 vss.t23 vss.t29 864.186
R137 vss.n80 vss.n79 855.515
R138 vss.n136 vss.n135 736.754
R139 vss.n51 vss.t23 655.605
R140 vss.n145 vss.n141 623.436
R141 vss.n143 vss.n141 623.436
R142 vss.n145 vss.n144 623.436
R143 vss.n144 vss.n143 623.436
R144 vss.n158 vss.n4 623.436
R145 vss.n160 vss.n4 623.436
R146 vss.n159 vss.n158 623.436
R147 vss.n160 vss.n159 623.436
R148 vss.n121 vss.n33 478.118
R149 vss.n135 vss.n134 451.765
R150 vss.n118 vss.n34 440.471
R151 vss.n163 vss.n162 421.781
R152 vss.n121 vss.n120 399.06
R153 vss.n136 vss.n9 399.034
R154 vss.n156 vss.t11 388.748
R155 vss.t17 vss.t9 378.079
R156 vss.n73 vss.n72 374.562
R157 vss.n150 vss.t36 373.755
R158 vss.t3 vss.t25 372.125
R159 vss.n113 vss.n40 356.894
R160 vss.n113 vss.n112 319.625
R161 vss.t3 vss.t7 309.608
R162 vss.t19 vss.t17 303.654
R163 vss.n92 vss.t19 302.166
R164 vss.t7 vss.n31 296.212
R165 vss.n69 vss.n48 292.5
R166 vss.n48 vss.t4 292.5
R167 vss.n49 vss.n47 292.5
R168 vss.n47 vss.t4 292.5
R169 vss.n76 vss.n45 292.5
R170 vss.n45 vss.t18 292.5
R171 vss.n46 vss.n44 292.5
R172 vss.n44 vss.t18 292.5
R173 vss.n112 vss.n39 292.5
R174 vss.n39 vss.t6 292.5
R175 vss.n40 vss.n38 292.5
R176 vss.n38 vss.t6 292.5
R177 vss.n153 vss.n150 292.5
R178 vss.n151 vss.n149 292.5
R179 vss.n149 vss.n148 292.5
R180 vss.n62 vss.n61 276.861
R181 vss.n61 vss.t25 233.695
R182 vss.t9 vss.n91 227.74
R183 vss.n89 vss.n85 219.482
R184 vss.n89 vss.n86 219.482
R185 vss.n94 vss.n86 219.482
R186 vss.n59 vss.n54 219.482
R187 vss.n56 vss.n54 219.482
R188 vss.n57 vss.n56 219.482
R189 vss.n116 vss.n37 215.702
R190 vss.n120 vss.n118 208.189
R191 vss.n56 vss.n55 195
R192 vss.n55 vss.n31 195
R193 vss.n60 vss.n59 195
R194 vss.n61 vss.n60 195
R195 vss.n94 vss.n93 195
R196 vss.n93 vss.n92 195
R197 vss.n90 vss.n89 195
R198 vss.n91 vss.n90 195
R199 vss.n92 vss.n37 165.083
R200 vss.t11 vss.n5 159.375
R201 vss.n58 vss.n57 134.776
R202 vss.n18 vss.n9 130.133
R203 vss.n95 vss.n85 128
R204 vss.n35 vss.n34 117.001
R205 vss.t0 vss.n35 117.001
R206 vss.n50 vss.n10 117.001
R207 vss.n51 vss.n50 117.001
R208 vss.n137 vss.n136 117.001
R209 vss.n138 vss.n137 117.001
R210 vss.n33 vss.n29 117.001
R211 vss.n62 vss.n29 117.001
R212 vss.n119 vss.n30 117.001
R213 vss.n37 vss.n30 117.001
R214 vss.n100 vss.n36 117.001
R215 vss.t0 vss.n36 117.001
R216 vss.n27 vss.n11 110.359
R217 vss.n115 vss.t6 107.85
R218 vss.n79 vss.t18 107.85
R219 vss.n73 vss.t18 107.85
R220 vss.n72 vss.t4 107.85
R221 vss.n66 vss.t4 107.85
R222 vss.n43 vss.t0 107.123
R223 vss.n95 vss.n94 91.4829
R224 vss.n107 vss.t1 86.2761
R225 vss.n106 vss.t33 86.2684
R226 vss.n16 vss.t24 86.2495
R227 vss.n23 vss.t26 85.2172
R228 vss.n96 vss.t20 85.2172
R229 vss.n91 vss.n32 84.8449
R230 vss.n80 vss.n43 80.1595
R231 vss.n116 vss.n115 78.7021
R232 vss.n59 vss.n58 78.0993
R233 vss.n21 vss.n11 73.4123
R234 vss.n128 vss.n24 68.9308
R235 vss.n14 vss.n13 68.8514
R236 vss.n63 vss.n62 68.4714
R237 vss.n106 vss.n105 68.1549
R238 vss.n16 vss.n15 68.0911
R239 vss.n14 vss.n12 68.0905
R240 vss.n65 vss.t36 65.8985
R241 vss.n83 vss.n40 65.3422
R242 vss.n147 vss.t28 58.5301
R243 vss.t28 vss.n5 58.5301
R244 vss.n156 vss.t36 58.5301
R245 vss.n162 vss.t36 58.5301
R246 vss.n57 vss.n53 58.5005
R247 vss.n53 vss.t3 58.5005
R248 vss.n54 vss.n52 58.5005
R249 vss.t3 vss.n52 58.5005
R250 vss.n88 vss.n85 58.5005
R251 vss.t17 vss.n88 58.5005
R252 vss.n87 vss.n86 58.5005
R253 vss.t17 vss.n87 58.5005
R254 vss.n100 vss.n82 55.9122
R255 vss.n161 vss.n160 48.7505
R256 vss.n162 vss.n161 48.7505
R257 vss.n158 vss.n157 48.7505
R258 vss.n157 vss.n156 48.7505
R259 vss.n143 vss.n142 48.7505
R260 vss.n142 vss.n5 48.7505
R261 vss.n146 vss.n145 48.7505
R262 vss.n147 vss.n146 48.7505
R263 vss.n111 vss.n110 45.5155
R264 vss.n123 vss.n31 44.6554
R265 vss.n102 vss.t12 44.1758
R266 vss.n103 vss.t5 43.3392
R267 vss.n125 vss.n28 33.5081
R268 vss.n111 vss.n41 30.4645
R269 vss.n123 vss.n32 28.282
R270 vss.n114 vss.n113 26.5914
R271 vss.n115 vss.n114 26.5914
R272 vss.n42 vss.n41 26.5914
R273 vss.n43 vss.n42 26.5914
R274 vss.n18 vss.n10 23.8938
R275 vss.n148 vss.n147 22.1468
R276 vss.n122 vss.n121 20.8934
R277 vss.n123 vss.n122 20.8934
R278 vss.n118 vss.n117 20.8934
R279 vss.n117 vss.n116 20.8934
R280 vss.n125 vss.n124 20.8934
R281 vss.n124 vss.n123 20.8934
R282 vss.n82 vss.n81 20.8934
R283 vss.n81 vss.n80 20.8934
R284 vss.n159 vss.n3 17.7278
R285 vss.n3 vss.t36 17.7278
R286 vss.n4 vss.n2 17.7278
R287 vss.n2 vss.t36 17.7278
R288 vss.n144 vss.n140 17.7278
R289 vss.n140 vss.t28 17.7278
R290 vss.n141 vss.n139 17.7278
R291 vss.n139 vss.t28 17.7278
R292 vss.n105 vss.t2 17.4005
R293 vss.n105 vss.t27 17.4005
R294 vss.n24 vss.t8 17.4005
R295 vss.n24 vss.t10 17.4005
R296 vss.n15 vss.t35 17.4005
R297 vss.n15 vss.t30 17.4005
R298 vss.n12 vss.t22 17.4005
R299 vss.n12 vss.t14 17.4005
R300 vss.n13 vss.t16 17.4005
R301 vss.n13 vss.t32 17.4005
R302 vss.n133 vss.n11 13.6763
R303 vss.n126 vss.n27 12.5161
R304 vss.n9 vss.n7 12.188
R305 vss.t13 vss.n7 12.188
R306 vss.n135 vss.n8 12.188
R307 vss.t13 vss.n8 12.188
R308 vss.n100 vss.n28 11.6757
R309 vss.n119 vss.n28 9.30959
R310 vss.n120 vss.n119 8.14595
R311 vss.n68 vss.n67 8.0142
R312 vss.n67 vss.n66 8.0142
R313 vss.n71 vss.n70 8.0142
R314 vss.n72 vss.n71 8.0142
R315 vss.n75 vss.n74 8.0142
R316 vss.n74 vss.n73 8.0142
R317 vss.n78 vss.n77 8.0142
R318 vss.n79 vss.n78 8.0142
R319 vss.n33 vss.n21 7.52991
R320 vss.n112 vss.n111 7.51354
R321 vss.n111 vss.n34 7.51354
R322 vss.n152 vss.n6 7.22272
R323 vss.t11 vss.n6 7.22272
R324 vss.n155 vss.n154 7.22272
R325 vss.t11 vss.n155 7.22272
R326 vss.n134 vss.n10 7.05622
R327 vss.n96 vss.n95 6.55702
R328 vss.n58 vss.n23 6.54313
R329 vss.n99 vss.n98 4.50397
R330 vss.n130 vss.n129 4.5005
R331 vss.n128 vss.n127 4.5005
R332 vss.n110 vss.n82 4.06119
R333 vss.n104 vss.n103 4.00099
R334 vss.n133 vss.n132 3.16116
R335 vss.n19 vss.n18 3.1005
R336 vss.n131 vss.n21 2.42272
R337 vss.n1 vss.n0 2.10264
R338 vss.n102 vss.n1 2.04087
R339 vss.n101 vss.n100 1.8605
R340 vss.n20 vss.n10 1.5505
R341 vss.n19 vss.n17 1.30682
R342 vss.n163 vss.n1 1.27326
R343 vss.n103 vss.n102 0.943777
R344 vss.n0 vss.t38 0.894893
R345 vss.t0 vss.t6 0.729218
R346 vss.n109 vss.n83 0.72262
R347 vss.n98 vss.n97 0.628972
R348 vss.n129 vss.n128 0.622028
R349 vss.n83 vss.n41 0.58329
R350 vss.n17 vss.n16 0.504667
R351 vss.n164 vss 0.441333
R352 vss.n108 vss.n104 0.379288
R353 vss.n110 vss.n109 0.358192
R354 vss.n127 vss.n126 0.344944
R355 vss.n129 vss.n23 0.311665
R356 vss.n98 vss.n96 0.308192
R357 vss vss.n164 0.274878
R358 vss.n17 vss.n14 0.263
R359 vss.n99 vss.n84 0.242521
R360 vss.n132 vss.n131 0.211936
R361 vss.n20 vss.n19 0.202941
R362 vss.n101 vss.n99 0.170929
R363 vss.n97 vss.n84 0.1505
R364 vss.n26 vss.n25 0.1505
R365 vss.n130 vss.n22 0.121511
R366 vss.n127 vss.n22 0.117521
R367 vss.n134 vss.n133 0.108289
R368 vss.n132 vss.n20 0.106883
R369 vss.n0 vss.t37 0.0927731
R370 vss.n27 vss.n22 0.0882358
R371 vss vss.n101 0.0866169
R372 vss.n108 vss.n107 0.0755
R373 vss.n131 vss.n130 0.063
R374 vss.n126 vss.n125 0.0573889
R375 vss vss.n163 0.0479585
R376 vss.n109 vss.n108 0.032697
R377 vss.n128 vss.n25 0.0143889
R378 vss.n104 vss 0.013548
R379 vss.n164 vss 0.0119108
R380 vss.n127 vss.n26 0.00581915
R381 vss.n107 vss.n106 0.00440625
R382 vss.n97 vss.n25 0.00397222
R383 vss.n84 vss.n26 0.00182979
R384 twin_tee_0.in.n2 twin_tee_0.in.t2 154.407
R385 twin_tee_0.in.n0 twin_tee_0.in.t0 43.1124
R386 twin_tee_0.in.n0 twin_tee_0.in.t1 10.2463
R387 twin_tee_0.in twin_tee_0.in.n5 9.43796
R388 twin_tee_0.in.n5 twin_tee_0.in.n4 4.5005
R389 twin_tee_0.in.n3 twin_tee_0.in.n1 2.2505
R390 twin_tee_0.in.n2 twin_tee_0.in.n1 1.48465
R391 twin_tee_0.in twin_tee_0.in.n0 0.723459
R392 twin_tee_0.in.n4 twin_tee_0.in.n2 0.394718
R393 twin_tee_0.in.n3 twin_tee_0.in 0.054875
R394 twin_tee_0.in.n5 twin_tee_0.in.n1 0.0307083
R395 twin_tee_0.in.n4 twin_tee_0.in.n3 0.002375
R396 twin_tee_0.c3_c4 twin_tee_0.c3_c4.t1 46.7014
R397 twin_tee_0.c3_c4 twin_tee_0.c3_c4.t0 0.349462
R398 twin_tee_0.c3_c4 twin_tee_0.c3_c4.n0 0.0354413
R399 twin_tee_0.c3_c4.n0 twin_tee_0.c3_c4.t2 0.0274722
R400 twin_tee_0.c3_c4.n0 twin_tee_0.c3_c4 0.0109069
R401 p3_opamp_0.VBIAS.n16 p3_opamp_0.VBIAS.n0 66.588
R402 p3_opamp_0.VBIAS.n13 p3_opamp_0.VBIAS.n1 66.588
R403 p3_opamp_0.VBIAS.n8 p3_opamp_0.VBIAS.t12 26.0899
R404 p3_opamp_0.VBIAS.n2 p3_opamp_0.VBIAS.t18 25.992
R405 p3_opamp_0.VBIAS.n7 p3_opamp_0.VBIAS.t13 25.5741
R406 p3_opamp_0.VBIAS.n11 p3_opamp_0.VBIAS.t7 25.5503
R407 p3_opamp_0.VBIAS.n14 p3_opamp_0.VBIAS.t5 25.5503
R408 p3_opamp_0.VBIAS.n15 p3_opamp_0.VBIAS.t3 25.5503
R409 p3_opamp_0.VBIAS.n17 p3_opamp_0.VBIAS.t1 25.5503
R410 p3_opamp_0.VBIAS.n2 p3_opamp_0.VBIAS.t16 25.5277
R411 p3_opamp_0.VBIAS.n3 p3_opamp_0.VBIAS.t14 25.5277
R412 p3_opamp_0.VBIAS.n4 p3_opamp_0.VBIAS.t19 25.5277
R413 p3_opamp_0.VBIAS.n5 p3_opamp_0.VBIAS.t17 25.5277
R414 p3_opamp_0.VBIAS.n6 p3_opamp_0.VBIAS.t15 25.5277
R415 p3_opamp_0.VBIAS.n8 p3_opamp_0.VBIAS.t9 25.5274
R416 p3_opamp_0.VBIAS.n9 p3_opamp_0.VBIAS.t10 25.5274
R417 p3_opamp_0.VBIAS.n10 p3_opamp_0.VBIAS.t11 25.5274
R418 p3_opamp_0.VBIAS.n0 p3_opamp_0.VBIAS.t2 17.4005
R419 p3_opamp_0.VBIAS.n0 p3_opamp_0.VBIAS.t4 17.4005
R420 p3_opamp_0.VBIAS.n1 p3_opamp_0.VBIAS.t6 17.4005
R421 p3_opamp_0.VBIAS.n1 p3_opamp_0.VBIAS.t8 17.4005
R422 p3_opamp_0.VBIAS.n12 p3_opamp_0.VBIAS.n7 7.30251
R423 p3_opamp_0.VBIAS p3_opamp_0.VBIAS.t0 3.31103
R424 p3_opamp_0.VBIAS.n11 p3_opamp_0.VBIAS.n10 1.19959
R425 p3_opamp_0.VBIAS.n10 p3_opamp_0.VBIAS.n9 0.6255
R426 p3_opamp_0.VBIAS.n9 p3_opamp_0.VBIAS.n8 0.583833
R427 p3_opamp_0.VBIAS.n3 p3_opamp_0.VBIAS.n2 0.5005
R428 p3_opamp_0.VBIAS.n5 p3_opamp_0.VBIAS.n4 0.482643
R429 p3_opamp_0.VBIAS.n6 p3_opamp_0.VBIAS.n5 0.464786
R430 p3_opamp_0.VBIAS.n4 p3_opamp_0.VBIAS.n3 0.429071
R431 p3_opamp_0.VBIAS p3_opamp_0.VBIAS.n17 0.197868
R432 p3_opamp_0.VBIAS.n15 p3_opamp_0.VBIAS.n14 0.151816
R433 p3_opamp_0.VBIAS.n7 p3_opamp_0.VBIAS.n6 0.136214
R434 p3_opamp_0.VBIAS.n14 p3_opamp_0.VBIAS.n13 0.0728684
R435 p3_opamp_0.VBIAS.n17 p3_opamp_0.VBIAS.n16 0.0728684
R436 p3_opamp_0.VBIAS.n16 p3_opamp_0.VBIAS.n15 0.0728684
R437 p3_opamp_0.VBIAS.n12 p3_opamp_0.VBIAS.n11 0.069579
R438 p3_opamp_0.VBIAS.n13 p3_opamp_0.VBIAS.n12 0.00378947
R439 p3_opamp_0.V1.n1 p3_opamp_0.V1.t8 240.631
R440 p3_opamp_0.V1.n0 p3_opamp_0.V1.t20 240.631
R441 p3_opamp_0.V1.n0 p3_opamp_0.V1.t7 240.349
R442 p3_opamp_0.V1.n0 p3_opamp_0.V1.t24 240.349
R443 p3_opamp_0.V1.n1 p3_opamp_0.V1.t16 240.349
R444 p3_opamp_0.V1.n1 p3_opamp_0.V1.t10 240.349
R445 p3_opamp_0.V1.n1 p3_opamp_0.V1.t12 240.349
R446 p3_opamp_0.V1.n1 p3_opamp_0.V1.t13 240.349
R447 p3_opamp_0.V1.n1 p3_opamp_0.V1.t9 240.349
R448 p3_opamp_0.V1.n1 p3_opamp_0.V1.t22 240.349
R449 p3_opamp_0.V1.n1 p3_opamp_0.V1.t14 240.349
R450 p3_opamp_0.V1.n0 p3_opamp_0.V1.t17 240.349
R451 p3_opamp_0.V1.n0 p3_opamp_0.V1.t21 240.349
R452 p3_opamp_0.V1.n0 p3_opamp_0.V1.t11 240.349
R453 p3_opamp_0.V1.n0 p3_opamp_0.V1.t25 240.349
R454 p3_opamp_0.V1.n0 p3_opamp_0.V1.t19 240.349
R455 p3_opamp_0.V1.n0 p3_opamp_0.V1.t23 240.349
R456 p3_opamp_0.V1.n0 p3_opamp_0.V1.t15 240.349
R457 p3_opamp_0.V1.n0 p3_opamp_0.V1.t18 240.349
R458 p3_opamp_0.V1.n0 p3_opamp_0.V1.t26 240.349
R459 p3_opamp_0.V1 p3_opamp_0.V1.t5 230.536
R460 p3_opamp_0.V1.n4 p3_opamp_0.V1.t4 229.337
R461 p3_opamp_0.V1 p3_opamp_0.V1.n3 201.905
R462 p3_opamp_0.V1 p3_opamp_0.V1.n2 201.904
R463 p3_opamp_0.V1.n4 p3_opamp_0.V1.t0 36.1494
R464 p3_opamp_0.V1.n3 p3_opamp_0.V1.t2 28.5655
R465 p3_opamp_0.V1.n3 p3_opamp_0.V1.t6 28.5655
R466 p3_opamp_0.V1.n2 p3_opamp_0.V1.t3 28.5655
R467 p3_opamp_0.V1.n2 p3_opamp_0.V1.t1 28.5655
R468 p3_opamp_0.V1 p3_opamp_0.V1.n0 8.1351
R469 p3_opamp_0.V1 p3_opamp_0.V1.n4 4.80549
R470 p3_opamp_0.V1.n0 p3_opamp_0.V1.n1 4.75675
R471 vdd.n50 vdd.n45 6857.65
R472 vdd.n50 vdd.n46 6857.65
R473 vdd.n48 vdd.n46 6857.65
R474 vdd.n48 vdd.n45 6857.65
R475 vdd.n11 vdd.n6 6130.59
R476 vdd.n11 vdd.n7 6130.59
R477 vdd.n9 vdd.n7 6130.59
R478 vdd.n9 vdd.n6 6130.59
R479 vdd.n25 vdd.n22 6130.59
R480 vdd.n25 vdd.n23 6130.59
R481 vdd.n27 vdd.n23 6130.59
R482 vdd.n27 vdd.n22 6130.59
R483 vdd.n47 vdd.n43 731.482
R484 vdd.n47 vdd.n44 731.482
R485 vdd.t60 vdd.t64 681.976
R486 vdd.t16 vdd.t60 681.976
R487 vdd.t12 vdd.t14 681.976
R488 vdd.t14 vdd.t8 681.976
R489 vdd.t2 vdd.t10 681.976
R490 vdd.t62 vdd.t2 681.976
R491 vdd.t4 vdd.t0 681.976
R492 vdd.t0 vdd.t6 681.976
R493 vdd.n8 vdd.n4 653.929
R494 vdd.n8 vdd.n5 653.929
R495 vdd.n24 vdd.n20 653.929
R496 vdd.n24 vdd.n21 653.929
R497 vdd.n51 vdd.n44 646.381
R498 vdd.n52 vdd.n43 625.601
R499 vdd.t64 vdd.n6 541.571
R500 vdd.t8 vdd.n7 541.571
R501 vdd.t10 vdd.n22 541.571
R502 vdd.t6 vdd.n23 541.571
R503 vdd.n12 vdd.n5 493.892
R504 vdd.n28 vdd.n21 487.142
R505 vdd.n13 vdd.n4 381.115
R506 vdd.n29 vdd.n20 372.925
R507 vdd.n10 vdd.t16 340.988
R508 vdd.n10 vdd.t12 340.988
R509 vdd.n26 vdd.t62 340.988
R510 vdd.n26 vdd.t4 340.988
R511 vdd.t55 vdd.n45 318.216
R512 vdd.t31 vdd.n46 318.216
R513 vdd.t39 vdd.t55 235.267
R514 vdd.t51 vdd.t39 235.267
R515 vdd.t47 vdd.t51 235.267
R516 vdd.t45 vdd.t47 235.267
R517 vdd.t53 vdd.t45 235.267
R518 vdd.t27 vdd.t53 235.267
R519 vdd.t43 vdd.t27 235.267
R520 vdd.t37 vdd.t43 235.267
R521 vdd.t29 vdd.t37 235.267
R522 vdd.t49 vdd.t21 235.267
R523 vdd.t21 vdd.t33 235.267
R524 vdd.t33 vdd.t25 235.267
R525 vdd.t25 vdd.t41 235.267
R526 vdd.t41 vdd.t35 235.267
R527 vdd.t35 vdd.t57 235.267
R528 vdd.t57 vdd.t23 235.267
R529 vdd.t23 vdd.t19 235.267
R530 vdd.t19 vdd.t31 235.267
R531 vdd.n34 vdd.t56 230.56
R532 vdd.n60 vdd.t32 230.405
R533 vdd.n15 vdd.n3 202.125
R534 vdd.n18 vdd.n1 201.834
R535 vdd.n16 vdd.n2 201.834
R536 vdd.n65 vdd.n56 201.779
R537 vdd.n35 vdd.n32 201.779
R538 vdd.n70 vdd.n41 201.761
R539 vdd.n34 vdd.n33 201.761
R540 vdd.n74 vdd.n37 201.761
R541 vdd.n73 vdd.n38 201.761
R542 vdd.n71 vdd.n40 201.761
R543 vdd.n66 vdd.n55 201.756
R544 vdd.n36 vdd.n31 201.756
R545 vdd.n63 vdd.n57 201.744
R546 vdd.n59 vdd.n58 201.744
R547 vdd.n72 vdd.n39 201.704
R548 vdd.n49 vdd.t29 117.633
R549 vdd.n49 vdd.t49 117.633
R550 vdd.n13 vdd.n12 44.5872
R551 vdd.n29 vdd.n28 43.1489
R552 vdd.n79 vdd.t59 43.0539
R553 vdd.n78 vdd.t18 42.7329
R554 vdd.n6 vdd.n4 30.8338
R555 vdd.n7 vdd.n5 30.8338
R556 vdd.n22 vdd.n20 30.8338
R557 vdd.n23 vdd.n21 30.8338
R558 vdd.n45 vdd.n43 30.8338
R559 vdd.n46 vdd.n44 30.8338
R560 vdd.n1 vdd.t65 28.5655
R561 vdd.n1 vdd.t61 28.5655
R562 vdd.n2 vdd.t17 28.5655
R563 vdd.n2 vdd.t13 28.5655
R564 vdd.n3 vdd.t15 28.5655
R565 vdd.n3 vdd.t9 28.5655
R566 vdd.n41 vdd.t22 28.5655
R567 vdd.n41 vdd.t34 28.5655
R568 vdd.n55 vdd.t26 28.5655
R569 vdd.n55 vdd.t42 28.5655
R570 vdd.n57 vdd.t36 28.5655
R571 vdd.n57 vdd.t58 28.5655
R572 vdd.n58 vdd.t24 28.5655
R573 vdd.n58 vdd.t20 28.5655
R574 vdd.n56 vdd.t1 28.5655
R575 vdd.n56 vdd.t7 28.5655
R576 vdd.n39 vdd.t63 28.5655
R577 vdd.n39 vdd.t5 28.5655
R578 vdd.n32 vdd.t11 28.5655
R579 vdd.n32 vdd.t3 28.5655
R580 vdd.n33 vdd.t40 28.5655
R581 vdd.n33 vdd.t52 28.5655
R582 vdd.n31 vdd.t48 28.5655
R583 vdd.n31 vdd.t46 28.5655
R584 vdd.n37 vdd.t54 28.5655
R585 vdd.n37 vdd.t28 28.5655
R586 vdd.n38 vdd.t44 28.5655
R587 vdd.n38 vdd.t38 28.5655
R588 vdd.n40 vdd.t30 28.5655
R589 vdd.n40 vdd.t50 28.5655
R590 vdd.n52 vdd.n51 15.3605
R591 vdd.n9 vdd.n8 4.5127
R592 vdd.n10 vdd.n9 4.5127
R593 vdd.n12 vdd.n11 4.5127
R594 vdd.n11 vdd.n10 4.5127
R595 vdd.n25 vdd.n24 4.5127
R596 vdd.n26 vdd.n25 4.5127
R597 vdd.n28 vdd.n27 4.5127
R598 vdd.n27 vdd.n26 4.5127
R599 vdd.n48 vdd.n47 3.85467
R600 vdd.n49 vdd.n48 3.85467
R601 vdd.n51 vdd.n50 3.85467
R602 vdd.n50 vdd.n49 3.85467
R603 vdd.n79 vdd 2.02508
R604 vdd.n67 vdd.n66 1.5005
R605 vdd.n70 vdd.n69 1.5005
R606 vdd.n61 vdd.n60 1.01532
R607 vdd.n19 vdd.n18 0.903037
R608 vdd.n77 vdd.n76 0.82517
R609 vdd.n68 vdd.n42 0.7505
R610 vdd.n64 vdd.n54 0.7505
R611 vdd vdd.n79 0.521599
R612 vdd.n18 vdd.n17 0.338735
R613 vdd.n17 vdd.n16 0.338735
R614 vdd.n14 vdd.n13 0.282318
R615 vdd.n30 vdd.n29 0.282318
R616 vdd.n15 vdd.n14 0.275967
R617 vdd.n16 vdd.n15 0.256696
R618 vdd.n74 vdd.n73 0.235794
R619 vdd.n71 vdd.n70 0.235794
R620 vdd.n53 vdd.n52 0.216779
R621 vdd.n75 vdd.n36 0.195353
R622 vdd.n77 vdd.n19 0.195317
R623 vdd.n60 vdd.n59 0.191472
R624 vdd.n63 vdd.n62 0.181056
R625 vdd.n19 vdd.n0 0.174399
R626 vdd.n17 vdd.n0 0.173577
R627 vdd.n62 vdd.n61 0.167167
R628 vdd.n61 vdd.n54 0.137765
R629 vdd.n35 vdd.n34 0.136529
R630 vdd.n78 vdd.n77 0.136138
R631 vdd.n72 vdd.n71 0.118147
R632 vdd.n64 vdd.n63 0.116513
R633 vdd.n70 vdd.n42 0.114471
R634 vdd.n66 vdd.n42 0.114471
R635 vdd.n73 vdd.n72 0.110794
R636 vdd.n69 vdd.n53 0.0996848
R637 vdd.n36 vdd.n35 0.0924118
R638 vdd.n66 vdd.n65 0.0924118
R639 vdd.n14 vdd.n0 0.0897857
R640 vdd.n76 vdd.n30 0.0888152
R641 vdd.n53 vdd.n30 0.0860978
R642 vdd.n76 vdd.n75 0.0755
R643 vdd vdd.n78 0.063
R644 vdd.n67 vdd.n54 0.0439783
R645 vdd.n69 vdd.n68 0.0426196
R646 vdd.n68 vdd.n67 0.0426196
R647 vdd.n62 vdd.n59 0.0421667
R648 vdd.n75 vdd.n74 0.0409412
R649 vdd.n65 vdd.n64 0.0262353
R650 p3_opamp_0.V2 p3_opamp_0.V2.t12 228.542
R651 p3_opamp_0.V2 p3_opamp_0.V2.t4 228.456
R652 p3_opamp_0.V2 p3_opamp_0.V2.n0 199.977
R653 p3_opamp_0.V2 p3_opamp_0.V2.n1 199.923
R654 p3_opamp_0.V2 p3_opamp_0.V2.t0 34.7182
R655 p3_opamp_0.V2.n0 p3_opamp_0.V2.t6 28.5655
R656 p3_opamp_0.V2.n0 p3_opamp_0.V2.t10 28.5655
R657 p3_opamp_0.V2.n1 p3_opamp_0.V2.t8 28.5655
R658 p3_opamp_0.V2.n1 p3_opamp_0.V2.t2 28.5655
R659 p3_opamp_0.V2 p3_opamp_0.V2.t3 26.6205
R660 p3_opamp_0.V2 p3_opamp_0.V2.t18 26.0942
R661 p3_opamp_0.V2 p3_opamp_0.V2.t14 26.0942
R662 p3_opamp_0.V2 p3_opamp_0.V2.t17 26.0942
R663 p3_opamp_0.V2 p3_opamp_0.V2.t16 26.0942
R664 p3_opamp_0.V2 p3_opamp_0.V2.t15 26.0942
R665 p3_opamp_0.V2 p3_opamp_0.V2.t13 26.0942
R666 p3_opamp_0.V2 p3_opamp_0.V2.t11 26.05
R667 p3_opamp_0.V2 p3_opamp_0.V2.t9 26.05
R668 p3_opamp_0.V2 p3_opamp_0.V2.t5 26.0489
R669 p3_opamp_0.V2 p3_opamp_0.V2.t1 26.0488
R670 p3_opamp_0.V2 p3_opamp_0.V2.t7 26.0478
C0 p3_opamp_0.VBIAS twin_tee_0.in 0.71001f
C1 out p3_opamp_0.VBIAS 2.97334f
C2 vdd p3_opamp_0.V2 14.0343f
C3 p3_opamp_0.PLUS p3_opamp_0.V2 0.04754f
C4 twin_tee_0.c3_c4 p3_opamp_0.V2 0.010504f
C5 p3_opamp_0.VX twin_tee_0.in 0.578867f
C6 out p3_opamp_0.VX 1.32e-21
C7 p3_opamp_0.V1 p3_opamp_0.V2 6.83344f
C8 p3_opamp_0.VX p3_opamp_0.VBIAS 1.88665f
C9 twin_tee_0.c3_c4 a_24144_17782# 0.257745f
C10 p3_opamp_0.PLUS vdd 0.52756f
C11 twin_tee_0.c3_c4 vdd 0.280465f
C12 p3_opamp_0.V2 twin_tee_0.in 0.55445f
C13 out p3_opamp_0.V2 0.004966f
C14 p3_opamp_0.V2 p3_opamp_0.VBIAS 0.190761f
C15 vdd p3_opamp_0.V1 9.40784f
C16 p3_opamp_0.PLUS p3_opamp_0.V1 0.654269f
C17 twin_tee_0.c3_c4 p3_opamp_0.V1 0.011866f
C18 p3_opamp_0.VX p3_opamp_0.V2 0.119464f
C19 a_24144_17782# twin_tee_0.in 1.64671f
C20 a_24144_17782# out 1.17749f
C21 vdd twin_tee_0.in 0.53616f
C22 p3_opamp_0.PLUS twin_tee_0.in 0.041f
C23 out vdd 5.12667f
C24 p3_opamp_0.PLUS out 0.455883f
C25 vdd p3_opamp_0.VBIAS 0.904256f
C26 p3_opamp_0.PLUS p3_opamp_0.VBIAS 0.738369f
C27 twin_tee_0.c3_c4 twin_tee_0.in 21.3079f
C28 twin_tee_0.c3_c4 out 21.970499f
C29 p3_opamp_0.V1 twin_tee_0.in 0.01158f
C30 out p3_opamp_0.V1 2.01513f
C31 p3_opamp_0.V1 p3_opamp_0.VBIAS 0.241132f
C32 p3_opamp_0.PLUS p3_opamp_0.VX 0.579422f
C33 p3_opamp_0.VX p3_opamp_0.V1 0.096512f
C34 out vss 16.742512f
C35 vdd vss 34.76173f
C36 p3_opamp_0.VX vss 1.45094f
C37 p3_opamp_0.V1 vss 12.79976f
C38 p3_opamp_0.V2 vss 21.56954f
C39 p3_opamp_0.VBIAS vss 26.706038f
C40 p3_opamp_0.PLUS vss 8.79069f
C41 twin_tee_0.c3_c4 vss 9.77697f
C42 twin_tee_0.in vss 21.124464f
C43 a_24144_17782# vss 57.9734f
C44 p3_opamp_0.V2.t0 vss 0.093093f
C45 p3_opamp_0.V2.t13 vss 0.456467f
C46 p3_opamp_0.V2.t12 vss 0.039293f
C47 p3_opamp_0.V2.t6 vss 0.01067f
C48 p3_opamp_0.V2.t10 vss 0.01067f
C49 p3_opamp_0.V2.n0 vss 0.022041f
C50 p3_opamp_0.V2.t8 vss 0.01067f
C51 p3_opamp_0.V2.t2 vss 0.01067f
C52 p3_opamp_0.V2.n1 vss 0.022034f
C53 p3_opamp_0.V2.t18 vss 0.456467f
C54 p3_opamp_0.V2.t14 vss 0.456467f
C55 p3_opamp_0.V2.t17 vss 0.456467f
C56 p3_opamp_0.V2.t16 vss 0.456467f
C57 p3_opamp_0.V2.t15 vss 0.456467f
C58 p3_opamp_0.V2.t4 vss 0.039293f
C59 p3_opamp_0.V2.t3 vss 0.45557f
C60 p3_opamp_0.V2.t7 vss 0.455564f
C61 p3_opamp_0.V2.t1 vss 0.45557f
C62 p3_opamp_0.V2.t5 vss 0.45557f
C63 p3_opamp_0.V2.t9 vss 0.45557f
C64 p3_opamp_0.V2.t11 vss 0.45557f
C65 vdd.t18 vss 0.019901f
C66 vdd.n0 vss 0.223596f
C67 vdd.t65 vss 0.005014f
C68 vdd.t61 vss 0.005014f
C69 vdd.n1 vss 0.010764f
C70 vdd.t17 vss 0.005014f
C71 vdd.t13 vss 0.005014f
C72 vdd.n2 vss 0.010764f
C73 vdd.t15 vss 0.005014f
C74 vdd.t9 vss 0.005014f
C75 vdd.n3 vss 0.011133f
C76 vdd.n4 vss 0.110301f
C77 vdd.n5 vss 0.105891f
C78 vdd.n6 vss 0.337331f
C79 vdd.n7 vss 0.337331f
C80 vdd.t64 vss 0.455865f
C81 vdd.t60 vss 0.505191f
C82 vdd.t16 vss 0.378893f
C83 vdd.t8 vss 0.455865f
C84 vdd.t14 vss 0.505191f
C85 vdd.t12 vss 0.378893f
C86 vdd.n8 vss 0.102411f
C87 vdd.n9 vss 0.102411f
C88 vdd.n10 vss 0.252596f
C89 vdd.n11 vss 0.102411f
C90 vdd.n12 vss 0.10405f
C91 vdd.n13 vss 0.096749f
C92 vdd.n14 vss 0.427321f
C93 vdd.n15 vss 0.676018f
C94 vdd.n16 vss 0.22694f
C95 vdd.n17 vss 0.1352f
C96 vdd.n18 vss 0.180024f
C97 vdd.n19 vss 0.310158f
C98 vdd.n20 vss 0.111125f
C99 vdd.n21 vss 0.10601f
C100 vdd.n22 vss 0.337331f
C101 vdd.n23 vss 0.337331f
C102 vdd.t10 vss 0.455865f
C103 vdd.t2 vss 0.505191f
C104 vdd.t62 vss 0.378893f
C105 vdd.n24 vss 0.102411f
C106 vdd.n25 vss 0.102411f
C107 vdd.t6 vss 0.455865f
C108 vdd.t0 vss 0.505191f
C109 vdd.t4 vss 0.378893f
C110 vdd.n26 vss 0.252596f
C111 vdd.n27 vss 0.102411f
C112 vdd.n28 vss 0.107685f
C113 vdd.n29 vss 0.100401f
C114 vdd.n30 vss 0.254494f
C115 vdd.t48 vss 0.005014f
C116 vdd.t46 vss 0.005014f
C117 vdd.n31 vss 0.010787f
C118 vdd.t11 vss 0.005014f
C119 vdd.t3 vss 0.005014f
C120 vdd.n32 vss 0.010772f
C121 vdd.t40 vss 0.005014f
C122 vdd.t52 vss 0.005014f
C123 vdd.n33 vss 0.010787f
C124 vdd.t56 vss 0.019032f
C125 vdd.n34 vss 0.348583f
C126 vdd.n35 vss 0.135105f
C127 vdd.n36 vss 0.158338f
C128 vdd.t54 vss 0.005014f
C129 vdd.t28 vss 0.005014f
C130 vdd.n37 vss 0.010787f
C131 vdd.t44 vss 0.005014f
C132 vdd.t38 vss 0.005014f
C133 vdd.n38 vss 0.010783f
C134 vdd.t63 vss 0.005014f
C135 vdd.t5 vss 0.005014f
C136 vdd.n39 vss 0.010759f
C137 vdd.t30 vss 0.005014f
C138 vdd.t50 vss 0.005014f
C139 vdd.n40 vss 0.010783f
C140 vdd.t22 vss 0.005014f
C141 vdd.t34 vss 0.005014f
C142 vdd.n41 vss 0.010787f
C143 vdd.n42 vss 0.045557f
C144 vdd.n43 vss 0.119518f
C145 vdd.n44 vss 0.120066f
C146 vdd.n45 vss 0.264865f
C147 vdd.n46 vss 0.264865f
C148 vdd.t55 vss 0.209561f
C149 vdd.t39 vss 0.17428f
C150 vdd.t51 vss 0.17428f
C151 vdd.t47 vss 0.17428f
C152 vdd.t45 vss 0.17428f
C153 vdd.t53 vss 0.17428f
C154 vdd.t27 vss 0.17428f
C155 vdd.t43 vss 0.17428f
C156 vdd.t37 vss 0.17428f
C157 vdd.t29 vss 0.13071f
C158 vdd.t31 vss 0.209561f
C159 vdd.t19 vss 0.17428f
C160 vdd.t23 vss 0.17428f
C161 vdd.t57 vss 0.17428f
C162 vdd.t35 vss 0.17428f
C163 vdd.t41 vss 0.17428f
C164 vdd.t25 vss 0.17428f
C165 vdd.t33 vss 0.17428f
C166 vdd.t21 vss 0.17428f
C167 vdd.t49 vss 0.13071f
C168 vdd.n47 vss 0.114488f
C169 vdd.n48 vss 0.114488f
C170 vdd.n49 vss 0.08714f
C171 vdd.n50 vss 0.114488f
C172 vdd.n51 vss 0.07041f
C173 vdd.n52 vss 0.068634f
C174 vdd.n53 vss 0.2704f
C175 vdd.n54 vss 0.21187f
C176 vdd.t26 vss 0.005014f
C177 vdd.t42 vss 0.005014f
C178 vdd.n55 vss 0.010787f
C179 vdd.t1 vss 0.005014f
C180 vdd.t7 vss 0.005014f
C181 vdd.n56 vss 0.010772f
C182 vdd.t36 vss 0.005014f
C183 vdd.t58 vss 0.005014f
C184 vdd.n57 vss 0.01078f
C185 vdd.t24 vss 0.005014f
C186 vdd.t20 vss 0.005014f
C187 vdd.n58 vss 0.010776f
C188 vdd.n59 vss 0.150396f
C189 vdd.t32 vss 0.018904f
C190 vdd.n60 vss 0.181286f
C191 vdd.n61 vss 0.35924f
C192 vdd.n62 vss 0.049792f
C193 vdd.n63 vss 0.164475f
C194 vdd.n64 vss 0.028491f
C195 vdd.n65 vss 0.113062f
C196 vdd.n66 vss 0.142172f
C197 vdd.n67 vss 0.125259f
C198 vdd.n68 vss 0.12327f
C199 vdd.n69 vss 0.206776f
C200 vdd.n70 vss 0.170828f
C201 vdd.n71 vss 0.170184f
C202 vdd.n72 vss 0.142725f
C203 vdd.n73 vss 0.168715f
C204 vdd.n74 vss 0.156133f
C205 vdd.n75 vss 0.047026f
C206 vdd.n76 vss 2.27976f
C207 vdd.n77 vss 2.04931f
C208 vdd.n78 vss 0.643573f
C209 vdd.t59 vss 0.021547f
C210 vdd.n79 vss 1.8034f
C211 p3_opamp_0.V1.n0 vss 1.40523f
C212 p3_opamp_0.V1.n1 vss 0.883305f
C213 p3_opamp_0.V1.t8 vss 0.215836f
C214 p3_opamp_0.V1.t16 vss 0.215719f
C215 p3_opamp_0.V1.t10 vss 0.215719f
C216 p3_opamp_0.V1.t12 vss 0.215719f
C217 p3_opamp_0.V1.t13 vss 0.215719f
C218 p3_opamp_0.V1.t9 vss 0.215719f
C219 p3_opamp_0.V1.t22 vss 0.215719f
C220 p3_opamp_0.V1.t14 vss 0.215719f
C221 p3_opamp_0.V1.t17 vss 0.215719f
C222 p3_opamp_0.V1.t21 vss 0.215719f
C223 p3_opamp_0.V1.t11 vss 0.215719f
C224 p3_opamp_0.V1.t25 vss 0.215719f
C225 p3_opamp_0.V1.t19 vss 0.215719f
C226 p3_opamp_0.V1.t23 vss 0.215719f
C227 p3_opamp_0.V1.t15 vss 0.215719f
C228 p3_opamp_0.V1.t18 vss 0.215719f
C229 p3_opamp_0.V1.t7 vss 0.215719f
C230 p3_opamp_0.V1.t20 vss 0.215838f
C231 p3_opamp_0.V1.t26 vss 0.215719f
C232 p3_opamp_0.V1.t24 vss 0.215719f
C233 p3_opamp_0.V1.t3 vss 0.017916f
C234 p3_opamp_0.V1.t1 vss 0.017916f
C235 p3_opamp_0.V1.n2 vss 0.038835f
C236 p3_opamp_0.V1.t2 vss 0.017916f
C237 p3_opamp_0.V1.t6 vss 0.017916f
C238 p3_opamp_0.V1.n3 vss 0.038818f
C239 p3_opamp_0.V1.t5 vss 0.069923f
C240 p3_opamp_0.V1.t0 vss 0.179078f
C241 p3_opamp_0.V1.t4 vss 0.066605f
C242 p3_opamp_0.V1.n4 vss 1.2521f
C243 p3_opamp_0.VBIAS.t0 vss 0.033592f
C244 p3_opamp_0.VBIAS.t2 vss 0.001609f
C245 p3_opamp_0.VBIAS.t4 vss 0.001609f
C246 p3_opamp_0.VBIAS.n0 vss 0.00353f
C247 p3_opamp_0.VBIAS.t6 vss 0.001609f
C248 p3_opamp_0.VBIAS.t8 vss 0.001609f
C249 p3_opamp_0.VBIAS.n1 vss 0.00353f
C250 p3_opamp_0.VBIAS.t18 vss 0.067433f
C251 p3_opamp_0.VBIAS.t16 vss 0.066149f
C252 p3_opamp_0.VBIAS.n2 vss 0.148179f
C253 p3_opamp_0.VBIAS.t14 vss 0.066149f
C254 p3_opamp_0.VBIAS.n3 vss 0.077179f
C255 p3_opamp_0.VBIAS.t19 vss 0.066149f
C256 p3_opamp_0.VBIAS.n4 vss 0.076984f
C257 p3_opamp_0.VBIAS.t17 vss 0.066149f
C258 p3_opamp_0.VBIAS.n5 vss 0.077373f
C259 p3_opamp_0.VBIAS.t15 vss 0.066149f
C260 p3_opamp_0.VBIAS.n6 vss 0.073605f
C261 p3_opamp_0.VBIAS.t13 vss 0.066286f
C262 p3_opamp_0.VBIAS.n7 vss 0.412165f
C263 p3_opamp_0.VBIAS.t12 vss 0.067681f
C264 p3_opamp_0.VBIAS.t9 vss 0.066142f
C265 p3_opamp_0.VBIAS.n8 vss 0.142758f
C266 p3_opamp_0.VBIAS.t10 vss 0.066142f
C267 p3_opamp_0.VBIAS.n9 vss 0.07339f
C268 p3_opamp_0.VBIAS.t11 vss 0.066142f
C269 p3_opamp_0.VBIAS.n10 vss 0.078801f
C270 p3_opamp_0.VBIAS.t7 vss 0.066241f
C271 p3_opamp_0.VBIAS.n11 vss 0.119554f
C272 p3_opamp_0.VBIAS.n12 vss 0.160208f
C273 p3_opamp_0.VBIAS.n13 vss 0.017329f
C274 p3_opamp_0.VBIAS.t5 vss 0.066241f
C275 p3_opamp_0.VBIAS.n14 vss 0.109887f
C276 p3_opamp_0.VBIAS.t3 vss 0.066241f
C277 p3_opamp_0.VBIAS.n15 vss 0.109887f
C278 p3_opamp_0.VBIAS.n16 vss 0.022864f
C279 p3_opamp_0.VBIAS.t1 vss 0.066241f
C280 p3_opamp_0.VBIAS.n17 vss 0.113577f
C281 twin_tee_0.c3_c4.t0 vss 14.727901f
C282 twin_tee_0.c3_c4.t2 vss 20.902302f
C283 twin_tee_0.c3_c4.n0 vss 6.25399f
C284 twin_tee_0.c3_c4.t1 vss 0.079662f
C285 twin_tee_0.in.t1 vss 16.2946f
C286 twin_tee_0.in.t0 vss 0.010986f
C287 twin_tee_0.in.n0 vss 0.979236f
C288 twin_tee_0.in.n1 vss 0.097937f
C289 twin_tee_0.in.t2 vss 0.045094f
C290 twin_tee_0.in.n2 vss 0.0445f
C291 twin_tee_0.in.n3 vss 0.008073f
C292 twin_tee_0.in.n4 vss 0.033356f
C293 twin_tee_0.in.n5 vss 1.40238f
C294 out.t1 vss 17.0627f
C295 out.t18 vss 0.030747f
C296 out.n0 vss 1.69316f
C297 out.n1 vss 0.319444f
C298 out.n2 vss 8.47466f
C299 out.n3 vss 0.228588f
C300 out.t23 vss 0.004354f
C301 out.t21 vss 0.004354f
C302 out.n4 vss 0.009991f
C303 out.t12 vss 0.004354f
C304 out.t4 vss 0.004354f
C305 out.n5 vss 0.009944f
C306 out.n6 vss 0.294111f
C307 out.t8 vss 0.015296f
C308 out.n7 vss 0.029896f
C309 out.t2 vss 0.004354f
C310 out.t9 vss 0.004354f
C311 out.n8 vss 0.009369f
C312 out.t13 vss 0.004354f
C313 out.t17 vss 0.004354f
C314 out.n9 vss 0.009307f
C315 out.t5 vss 0.004354f
C316 out.t10 vss 0.004354f
C317 out.n10 vss 0.009296f
C318 out.t22 vss 0.004354f
C319 out.t14 vss 0.004354f
C320 out.n11 vss 0.010391f
C321 out.t25 vss 0.004354f
C322 out.t16 vss 0.004354f
C323 out.n12 vss 0.009296f
C324 out.t3 vss 0.004354f
C325 out.t20 vss 0.004354f
C326 out.n13 vss 0.009296f
C327 out.t6 vss 0.004354f
C328 out.t24 vss 0.004354f
C329 out.n14 vss 0.009296f
C330 out.t7 vss 0.004354f
C331 out.t27 vss 0.004354f
C332 out.n15 vss 0.010471f
C333 out.t0 vss 0.004354f
C334 out.t28 vss 0.004354f
C335 out.n16 vss 0.009288f
C336 out.t26 vss 0.004354f
C337 out.t11 vss 0.004354f
C338 out.n17 vss 0.009288f
C339 out.t19 vss 0.004354f
C340 out.t15 vss 0.004354f
C341 out.n18 vss 0.011309f
C342 out.n19 vss 0.411658f
C343 out.n20 vss 0.143381f
C344 out.n21 vss 0.157433f
C345 out.n22 vss 0.179935f
C346 out.n23 vss 0.189695f
C347 out.n24 vss 0.915709f
C348 out.n25 vss 0.155485f
C349 out.n26 vss 0.184815f
C350 out.n27 vss 0.173542f
C351 out.n28 vss 0.143412f
C352 out.n29 vss 0.722411f
C353 out.n30 vss 0.351424f
C354 out.n31 vss 3.85203f
.ends

