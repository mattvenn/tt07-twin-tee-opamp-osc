VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO twin_tee
  CLASS BLOCK ;
  FOREIGN twin_tee ;
  ORIGIN 3.840 19.190 ;
  SIZE 45.140 BY 46.360 ;
  PIN vss
    ANTENNADIFFAREA 6.709700 ;
    PORT
      LAYER met1 ;
        RECT -3.080 14.300 -2.080 15.300 ;
    END
  END vss
  PIN out
    PORT
      LAYER met1 ;
        RECT 39.510 25.020 40.510 26.020 ;
    END
  END out
  PIN in
    PORT
      LAYER met1 ;
        RECT -3.130 25.060 -2.130 26.060 ;
    END
  END in
  OBS
      LAYER pwell ;
        RECT 3.660 20.890 16.120 26.220 ;
        RECT 22.450 20.950 34.910 26.280 ;
        RECT 6.280 -19.190 35.260 -17.180 ;
      LAYER li1 ;
        RECT 3.840 25.870 15.940 26.040 ;
        RECT 3.840 21.240 4.010 25.870 ;
        RECT 4.840 25.390 7.190 25.450 ;
        RECT 4.490 25.040 7.190 25.390 ;
        RECT 4.840 24.940 7.190 25.040 ;
        RECT 12.690 22.070 15.050 22.110 ;
        RECT 12.690 21.720 15.290 22.070 ;
        RECT 12.690 21.600 15.050 21.720 ;
        RECT 15.770 21.240 15.940 25.870 ;
        RECT 3.840 21.070 15.940 21.240 ;
        RECT 22.630 25.930 34.730 26.100 ;
        RECT 22.630 21.300 22.800 25.930 ;
        RECT 23.520 25.450 25.880 25.540 ;
        RECT 23.280 25.100 25.880 25.450 ;
        RECT 23.520 25.020 25.880 25.100 ;
        RECT 31.340 22.130 33.730 22.230 ;
        RECT 31.340 21.780 34.080 22.130 ;
        RECT 31.340 21.710 33.730 21.780 ;
        RECT 34.560 21.300 34.730 25.930 ;
        RECT 22.630 21.130 34.730 21.300 ;
        RECT -2.280 16.500 0.010 19.350 ;
        RECT 6.460 -17.530 35.080 -17.360 ;
        RECT 6.460 -18.840 6.630 -17.530 ;
        RECT 7.050 -18.390 9.290 -17.920 ;
        RECT 32.230 -18.390 34.460 -17.950 ;
        RECT 34.910 -18.840 35.080 -17.530 ;
        RECT 6.460 -19.010 35.080 -18.840 ;
      LAYER mcon ;
        RECT -2.280 16.880 0.010 18.870 ;
      LAYER met1 ;
        RECT -3.840 26.060 -1.570 26.490 ;
        RECT -3.840 25.060 -3.130 26.060 ;
        RECT -2.130 25.580 -1.570 26.060 ;
        RECT 39.030 26.020 41.300 27.170 ;
        RECT 39.030 25.815 39.510 26.020 ;
        RECT -2.130 25.060 7.300 25.580 ;
        RECT -3.840 24.840 7.300 25.060 ;
        RECT 17.250 24.930 26.180 25.610 ;
        RECT 36.615 25.185 39.510 25.815 ;
        RECT -3.840 23.980 -1.570 24.840 ;
        RECT 1.880 19.690 2.620 24.840 ;
        RECT 17.250 22.180 17.930 24.930 ;
        RECT 36.615 22.290 37.245 25.185 ;
        RECT 38.890 25.020 39.510 25.185 ;
        RECT 40.510 25.020 41.300 26.020 ;
        RECT 38.890 24.660 41.300 25.020 ;
        RECT 12.520 21.500 19.540 22.180 ;
        RECT 31.270 21.660 37.270 22.290 ;
        RECT 38.890 19.760 39.835 24.660 ;
        RECT -2.430 16.210 0.210 19.270 ;
        RECT 1.880 18.950 9.940 19.690 ;
        RECT -3.300 15.300 0.210 16.210 ;
        RECT -3.300 14.300 -3.080 15.300 ;
        RECT -2.080 14.300 0.210 15.300 ;
        RECT -3.300 13.800 0.210 14.300 ;
        RECT -3.300 13.700 -1.030 13.800 ;
        RECT -2.810 2.045 -1.620 13.700 ;
        RECT -2.810 0.855 4.705 2.045 ;
        RECT -2.810 -17.780 -1.620 0.855 ;
        RECT -1.080 0.850 2.000 0.855 ;
        RECT 9.210 0.530 9.930 18.950 ;
        RECT 38.810 15.920 39.910 19.760 ;
        RECT 38.780 14.820 39.940 15.920 ;
        RECT 4.180 -0.190 9.930 0.530 ;
        RECT 19.110 -15.920 19.890 -10.570 ;
        RECT 19.110 -16.700 37.650 -15.920 ;
        RECT -2.810 -18.535 9.415 -17.780 ;
        RECT 36.870 -17.820 37.650 -16.700 ;
        RECT -2.810 -18.755 -1.620 -18.535 ;
        RECT 32.100 -18.600 37.650 -17.820 ;
      LAYER via ;
        RECT 18.830 21.500 19.510 22.180 ;
        RECT 3.485 0.855 4.675 2.045 ;
        RECT 38.810 14.820 39.910 15.920 ;
        RECT 4.210 -0.190 4.930 0.530 ;
        RECT 19.110 -11.380 19.890 -10.600 ;
      LAYER met2 ;
        RECT 18.830 20.375 19.510 22.210 ;
        RECT 38.810 12.405 39.910 15.950 ;
        RECT 38.790 11.355 39.930 12.405 ;
        RECT 38.810 11.330 39.910 11.355 ;
        RECT 3.485 2.045 4.675 2.075 ;
        RECT 3.485 0.855 6.560 2.045 ;
        RECT 3.485 0.825 4.675 0.855 ;
        RECT 4.210 0.530 4.930 0.560 ;
        RECT 0.385 -0.190 4.930 0.530 ;
        RECT 4.210 -0.220 4.930 -0.190 ;
        RECT 19.110 -10.600 19.890 -8.555 ;
        RECT 19.080 -11.380 19.920 -10.600 ;
      LAYER via2 ;
        RECT 18.830 20.420 19.510 21.100 ;
        RECT 38.835 11.355 39.885 12.405 ;
        RECT 5.325 0.855 6.515 2.045 ;
        RECT 0.430 -0.190 1.150 0.530 ;
        RECT 19.110 -9.380 19.890 -8.600 ;
      LAYER met3 ;
        RECT 18.805 20.395 19.535 21.125 ;
        RECT 18.830 19.600 19.510 20.395 ;
        RECT 1.745 2.735 18.605 18.135 ;
        RECT 20.490 2.550 37.350 17.950 ;
        RECT 5.300 2.045 6.540 2.070 ;
        RECT 5.300 0.855 8.085 2.045 ;
        RECT 5.300 0.830 6.540 0.855 ;
        RECT 38.810 0.795 39.910 12.430 ;
        RECT 0.405 -0.215 1.175 0.555 ;
        RECT 0.430 -2.350 1.150 -0.215 ;
        RECT 1.700 -15.860 18.560 -0.460 ;
        RECT 19.110 -8.575 19.890 -6.980 ;
        RECT 19.085 -9.405 19.915 -8.575 ;
        RECT 20.660 -15.660 37.520 -0.260 ;
        RECT 38.785 -0.295 39.935 0.795 ;
        RECT 38.810 -0.300 39.910 -0.295 ;
      LAYER via3 ;
        RECT 18.830 19.630 19.510 20.310 ;
        RECT 18.185 2.875 18.505 17.995 ;
        RECT 36.930 2.690 37.250 17.810 ;
        RECT 6.865 0.855 8.055 2.045 ;
        RECT 38.815 -0.295 39.905 0.795 ;
        RECT 0.430 -2.320 1.150 -1.600 ;
        RECT 18.140 -15.720 18.460 -0.600 ;
        RECT 19.110 -7.790 19.890 -7.010 ;
        RECT 37.100 -15.520 37.420 -0.400 ;
      LAYER met4 ;
        RECT 18.825 19.820 19.515 20.315 ;
        RECT 17.710 18.640 37.680 19.820 ;
        RECT 2.140 3.130 16.750 17.740 ;
        RECT 17.710 12.800 18.890 18.640 ;
        RECT 8.580 2.085 9.710 3.130 ;
        RECT 18.105 2.795 18.585 12.800 ;
        RECT 20.885 2.945 35.495 17.555 ;
        RECT 36.500 12.240 37.680 18.640 ;
        RECT 28.575 2.085 29.705 2.945 ;
        RECT 36.850 2.610 37.330 12.240 ;
        RECT 6.860 2.045 8.060 2.050 ;
        RECT 8.580 2.045 29.705 2.085 ;
        RECT 6.860 0.955 29.705 2.045 ;
        RECT 6.860 0.855 9.505 0.955 ;
        RECT 6.860 0.850 8.060 0.855 ;
        RECT 36.670 -0.300 39.910 0.800 ;
        RECT 0.425 -2.325 1.155 -1.595 ;
        RECT 0.430 -2.850 1.150 -2.325 ;
        RECT 2.095 -2.850 16.705 -0.855 ;
        RECT 18.060 -0.980 18.540 -0.520 ;
        RECT 21.055 -0.980 35.665 -0.655 ;
        RECT 0.430 -3.570 16.705 -2.850 ;
        RECT 2.095 -15.465 16.705 -3.570 ;
        RECT 17.820 -5.790 35.665 -0.980 ;
        RECT 36.670 -5.140 37.770 -0.300 ;
        RECT 18.060 -15.800 18.540 -5.790 ;
        RECT 19.110 -7.005 19.890 -5.790 ;
        RECT 19.105 -7.795 19.895 -7.005 ;
        RECT 21.055 -15.265 35.665 -5.790 ;
        RECT 37.020 -15.600 37.500 -5.140 ;
  END
END twin_tee
END LIBRARY

